// RUN: eqmap %s -f -t 8 %s.opt && equiv_fpga %s.opt %s | FileCheck %s && rm %s.opt

// Verilog
// c7552
// Ninputs 207
// Noutputs 108
// NtotalGates 3513
// BUFF1 535
// NOT1 876
// AND2 534
// AND4 64
// NAND2 1028
// NOR2 40
// OR2 180
// OR3 10
// AND5 32
// AND3 146
// OR5 24
// OR4 30
// NOR3 10
// NOR4 4

// CHECK: Equivalence successfully proven!

module c7552 (
    N1,
    N5,
    N9,
    N12,
    N15,
    N18,
    N23,
    N26,
    N29,
    N32,
    N35,
    N38,
    N41,
    N44,
    N47,
    N50,
    N53,
    N54,
    N55,
    N56,
    N57,
    N58,
    N59,
    N60,
    N61,
    N62,
    N63,
    N64,
    N65,
    N66,
    N69,
    N70,
    N73,
    N74,
    N75,
    N76,
    N77,
    N78,
    N79,
    N80,
    N81,
    N82,
    N83,
    N84,
    N85,
    N86,
    N87,
    N88,
    N89,
    N94,
    N97,
    N100,
    N103,
    N106,
    N109,
    N110,
    N111,
    N112,
    N113,
    N114,
    N115,
    N118,
    N121,
    N124,
    N127,
    N130,
    N133,
    N134,
    N135,
    N138,
    N141,
    N144,
    N147,
    N150,
    N151,
    N152,
    N153,
    N154,
    N155,
    N156,
    N157,
    N158,
    N159,
    N160,
    N161,
    N162,
    N163,
    N164,
    N165,
    N166,
    N167,
    N168,
    N169,
    N170,
    N171,
    N172,
    N173,
    N174,
    N175,
    N176,
    N177,
    N178,
    N179,
    N180,
    N181,
    N182,
    N183,
    N184,
    N185,
    N186,
    N187,
    N188,
    N189,
    N190,
    N191,
    N192,
    N193,
    N194,
    N195,
    N196,
    N197,
    N198,
    N199,
    N200,
    N201,
    N202,
    N203,
    N204,
    N205,
    N206,
    N207,
    N208,
    N209,
    N210,
    N211,
    N212,
    N213,
    N214,
    N215,
    N216,
    N217,
    N218,
    N219,
    N220,
    N221,
    N222,
    N223,
    N224,
    N225,
    N226,
    N227,
    N228,
    N229,
    N230,
    N231,
    N232,
    N233,
    N234,
    N235,
    N236,
    N237,
    N238,
    N239,
    N240,
    N242,
    N245,
    N248,
    N251,
    N254,
    N257,
    N260,
    N263,
    N267,
    N271,
    N274,
    N277,
    N280,
    N283,
    N286,
    N289,
    N293,
    N296,
    N299,
    N303,
    N307,
    N310,
    N313,
    N316,
    N319,
    N322,
    N325,
    N328,
    N331,
    N334,
    N337,
    N340,
    N343,
    N346,
    N349,
    N352,
    N355,
    N358,
    N361,
    N364,
    N367,
    N382,
    N241_I,
    N387,
    N388,
    N478,
    N482,
    N484,
    N486,
    N489,
    N492,
    N501,
    N505,
    N507,
    N509,
    N511,
    N513,
    N515,
    N517,
    N519,
    N535,
    N537,
    N539,
    N541,
    N543,
    N545,
    N547,
    N549,
    N551,
    N553,
    N556,
    N559,
    N561,
    N563,
    N565,
    N567,
    N569,
    N571,
    N573,
    N582,
    N643,
    N707,
    N813,
    N881,
    N882,
    N883,
    N884,
    N885,
    N889,
    N945,
    N1110,
    N1111,
    N1112,
    N1113,
    N1114,
    N1489,
    N1490,
    N1781,
    N10025,
    N10101,
    N10102,
    N10103,
    N10104,
    N10109,
    N10110,
    N10111,
    N10112,
    N10350,
    N10351,
    N10352,
    N10353,
    N10574,
    N10575,
    N10576,
    N10628,
    N10632,
    N10641,
    N10704,
    N10706,
    N10711,
    N10712,
    N10713,
    N10714,
    N10715,
    N10716,
    N10717,
    N10718,
    N10729,
    N10759,
    N10760,
    N10761,
    N10762,
    N10763,
    N10827,
    N10837,
    N10838,
    N10839,
    N10840,
    N10868,
    N10869,
    N10870,
    N10871,
    N10905,
    N10906,
    N10907,
    N10908,
    N11333,
    N11334,
    N11340,
    N11342,
    N241_O
);

  input N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
      N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
      N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
      N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
      N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
      N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
      N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
      N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
      N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
      N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
      N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
      N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
      N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
      N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
      N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
      N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
      N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
      N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
      N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
      N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
      N355,N358,N361,N364,N367,N382,N241_I;

  output N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,
       N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,
       N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,
       N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,
       N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,
       N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,
       N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,
       N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,
       N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,
       N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,
       N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O;

  wire N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,
     N599,N604,N609,N614,N625,N628,N632,N636,N641,N642,
     N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,
     N688,N689,N695,N700,N705,N706,N708,N715,N721,N727,
     N733,N734,N742,N748,N749,N750,N758,N759,N762,N768,
     N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,
     N833,N839,N845,N853,N859,N865,N871,N886,N887,N957,
     N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,
     N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,
     N1206,N1211,N1218,N1222,N1227,N1233,N1240,N1244,N1249,N1256,
     N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,
     N1305,N1308,N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,
     N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,N1359,N1362,
     N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,
     N1395,N1398,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,
     N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,
     N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,
     N1485,N1537,N1551,N1649,N1703,N1708,N1713,N1721,N1758,N1782,
     N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,
     N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,
     N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,N1835,N1839,
     N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,
     N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,
     N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
     N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,
     N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,
     N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,
     N1946,N1947,N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,
     N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
     N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,
     N1995,N1996,N1997,N2003,N2010,N2011,N2012,N2013,N2014,N2015,
     N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,
     N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,
     N2070,N2071,N2072,N2073,N2074,N2081,N2086,N2107,N2108,N2110,
     N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,
     N2235,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
     N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,
     N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,
     N2282,N2283,N2284,N2285,N2286,N2287,N2293,N2299,N2300,N2301,
     N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,
     N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,
     N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,
     N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,
     N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
     N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,
     N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,
     N2402,N2403,N2404,N2405,N2406,N2412,N2418,N2419,N2420,N2421,
     N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
     N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,
     N2454,N2458,N2462,N2466,N2470,N2474,N2478,N2482,N2488,N2496,
     N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,
     N2561,N2567,N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,
     N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,N2670,N2674,
     N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,
     N2741,N2745,N2749,N2753,N2757,N2761,N2765,N2766,N2769,N2772,
     N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,
     N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,
     N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,
     N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,
     N3006,N3007,N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,
     N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,N3036,N3037,
     N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,
     N3096,N3097,N3101,N3107,N3114,N3122,N3126,N3130,N3131,N3134,
     N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,
     N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,
     N3215,N3221,N3228,N3229,N3232,N3236,N3241,N3247,N3251,N3255,
     N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,
     N3311,N3315,N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,
     N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,
     N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,
     N3404,N3410,N3416,N3420,N3424,N3428,N3432,N3436,N3440,N3444,
     N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,
     N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,
     N3515,N3518,N3521,N3524,N3527,N3530,N3535,N3539,N3542,N3545,
     N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,
     N3571,N3574,N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,
     N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,N3625,N3628,
     N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,
     N3661,N3664,N3667,N3670,N3673,N3676,N3679,N3682,N3685,N3688,
     N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,
     N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,
     N3751,N3754,N3757,N3760,N3763,N3766,N3769,N3772,N3775,N3778,
     N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,
     N3807,N3810,N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,
     N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,N3861,N3864,
     N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,
     N3954,N3955,N3956,N3958,N3964,N4193,N4303,N4308,N4313,N4326,
     N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,
     N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
     N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,
     N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,
     N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,
     N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
     N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,
     N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,
     N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,
     N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,
     N4593,N4597,N4603,N4610,N4611,N4612,N4613,N4614,N4615,N4616,
     N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,
     N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,
     N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,
     N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,
     N4667,N4674,N4675,N4678,N4682,N4687,N4693,N4694,N4695,N4696,
     N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,
     N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,
     N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,
     N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,
     N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
     N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,N4801,N4802,
     N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,
     N4829,N4832,N4835,N4838,N4841,N4844,N4847,N4850,N4853,N4856,
     N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,
     N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,
     N4919,N4922,N4925,N4928,N4931,N4934,N4937,N4940,N4943,N4946,
     N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,
     N4979,N4982,N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,
     N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,N5033,N5036,
     N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,
     N5061,N5064,N5065,N5066,N5067,N5068,N5071,N5074,N5077,N5080,
     N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,
     N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,
     N5135,N5138,N5141,N5144,N5147,N5150,N5153,N5156,N5159,N5162,
     N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,
     N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
     N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5196,
     N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,
     N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5283,N5284,N5285,
     N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,
     N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,
     N5319,N5320,N5321,N5322,N5323,N5324,N5363,N5364,N5365,N5366,
     N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,
     N5452,N5453,N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,
     N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,N5587,N5602,
     N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,
     N5697,N5707,N5718,N5728,N5735,N5736,N5740,N5744,N5747,N5751,
     N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,
     N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,
     N5905,N5915,N5926,N5936,N5943,N5944,N5945,N5946,N5947,N5948,
     N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,
     N5959,N5960,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,
     N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5989,N5990,
     N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,
     N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,
     N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,
     N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,
     N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
     N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,
     N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,
     N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,
     N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,
     N6126,N6127,N6131,N6135,N6136,N6137,N6141,N6145,N6148,N6149,
     N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,
     N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,
     N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,
     N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,
     N6207,N6210,N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,
     N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,N6239,N6240,
     N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,
     N6259,N6260,N6261,N6262,N6263,N6266,N6540,N6541,N6542,N6543,
     N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,
     N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,
     N6602,N6603,N6604,N6605,N6606,N6621,N6622,N6623,N6624,N6625,
     N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,
     N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,
     N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,N6677,N6678,
     N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,
     N6689,N6690,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,
     N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,
     N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,
     N6756,N6757,N6758,N6761,N6762,N6766,N6767,N6768,N6769,N6770,
     N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,
     N6781,N6782,N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,
     N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,N6809,N6812,
     N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,
     N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6848,N6849,N6850,
     N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,
     N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,
     N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6884,
     N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,
     N6901,N6912,N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,
     N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,N7055,N7056,
     N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
     N7073,N7077,N7080,N7086,N7091,N7095,N7098,N7099,N7100,N7103,
     N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,
     N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,
     N7213,N7216,N7219,N7222,N7229,N7240,N7250,N7258,N7272,N7288,
     N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,
     N7340,N7343,N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,
     N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,N7402,N7405,
     N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,
     N7438,N7441,N7444,N7447,N7450,N7453,N7456,N7459,N7462,N7465,
     N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,
     N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,
     N7524,N7527,N7530,N7533,N7536,N7539,N7542,N7545,N7548,N7551,
     N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,
     N7572,N7573,N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,
     N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,N7671,N7744,
     N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,
     N8146,N8156,N8166,N8169,N8183,N8186,N8196,N8200,N8204,N8208,
     N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,
     N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,
     N8261,N8262,N8269,N8274,N8275,N8276,N8277,N8278,N8279,N8280,
     N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,
     N8298,N8307,N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,
     N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,
     N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,
     N8355,N8356,N8357,N8358,N8365,N8369,N8370,N8371,N8372,N8373,
     N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,
     N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,
     N8394,N8404,N8405,N8409,N8410,N8411,N8412,N8415,N8416,N8417,
     N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,
     N8440,N8441,N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,
     N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,N8466,N8469,
     N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,
     N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8500,N8501,
     N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,
     N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,
     N8528,N8531,N8534,N8537,N8538,N8539,N8540,N8541,N8545,N8546,
     N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,
     N8565,N8566,N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,
     N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,N8609,N8610,
     N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,
     N8633,N8634,N8637,N8638,N8639,N8644,N8645,N8646,N8647,N8648,
     N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,
     N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,
     N8711,N8714,N8717,N8718,N8721,N8724,N8727,N8730,N8733,N8734,
     N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,
     N8757,N8760,N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,
     N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,N8811,N8814,
     N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,
     N8865,N8866,N8871,N8874,N8878,N8879,N8880,N8881,N8882,N8883,
     N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,
     N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,
     N8995,N8996,N9001,N9005,N9024,N9025,N9029,N9035,N9053,N9054,
     N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,
     N9079,N9082,N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,
     N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,N9146,N9149,
     N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,
     N9183,N9193,N9203,N9206,N9220,N9223,N9234,N9235,N9236,N9237,
     N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,
     N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,
     N9268,N9271,N9272,N9273,N9274,N9275,N9276,N9280,N9285,N9286,
     N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,
     N9301,N9307,N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,
     N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,N9358,N9359,
     N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,
     N9370,N9371,N9372,N9375,N9381,N9382,N9383,N9384,N9385,N9392,
     N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,
     N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,
     N9420,N9421,N9422,N9423,N9426,N9429,N9432,N9435,N9442,N9445,
     N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,
     N9468,N9473,N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,
     N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,N9514,N9515,
     N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,
     N9555,N9556,N9557,N9560,N9561,N9562,N9563,N9564,N9565,N9566,
     N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,
     N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,
     N9601,N9602,N9603,N9604,N9605,N9608,N9611,N9612,N9613,N9614,
     N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,
     N9632,N9635,N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,
     N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,N9674,N9675,
     N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,
     N9707,N9710,N9711,N9714,N9715,N9716,N9717,N9720,N9721,N9722,
     N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
     N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,
     N9766,N9767,N9768,N9769,N9773,N9774,N9775,N9779,N9784,N9785,
     N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,
     N9802,N9803,N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,
     N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,N9836,N9837,
     N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,
     N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,
     N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,
     N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,
     N9947,N9948,N9949,N9953,N9954,N9955,N9956,N9957,N9958,N9959,
     N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,
     N9974,N9975,N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,
     N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,N10006,N10007,
     N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,
     N10022,N10023,N10024,N10026,N10028,N10032,N10033,N10034,N10035,N10036,
     N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,
     N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,
     N10073,N10076,N10077,N10082,N10083,N10084,N10085,N10086,N10093,N10094,
     N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,
     N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,
     N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,N10160,N10161,
     N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,
     N10180,N10183,N10186,N10189,N10192,N10195,N10196,N10197,N10200,N10203,
     N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,
     N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,
     N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10278,
     N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,
     N10292,N10293,N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,
     N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,N10324,N10325,
     N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,
     N10338,N10339,N10340,N10341,N10344,N10354,N10357,N10360,N10367,N10375,
     N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,
     N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,
     N10444,N10445,N10450,N10451,N10455,N10456,N10465,N10466,N10479,N10497,
     N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,
     N10531,N10534,N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,
     N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,
     N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,
     N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10577,N10581,N10582,
     N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,
     N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,
     N10640,N10642,N10643,N10644,N10645,N10647,N10648,N10649,N10652,N10659,
     N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,
     N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,
     N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,N10708,N10709,
     N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,
     N10748,N10749,N10750,N10753,N10754,N10764,N10765,N10766,N10767,N10768,
     N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,
     N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,
     N10809,N10812,N10815,N10816,N10817,N10820,N10823,N10824,N10825,N10826,
     N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,
     N10864,N10865,N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,
     N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,N10890,N10891,
     N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,
     N10916,N10917,N10918,N10919,N10922,N10923,N10928,N10931,N10934,N10935,
     N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,
     N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,
     N10988,N10989,N10990,N10991,N10992,N10995,N10998,N10999,N11000,N11001,
     N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,
     N11014,N11015,N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,
     N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,N11050,N11053,
     N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,
     N11076,N11077,N11078,N11095,N11098,N11099,N11100,N11103,N11106,N11107,
     N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,
     N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,
     N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11152,N11153,
     N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,
     N11180,N11183,N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,
     N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,N11222,
     N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,
     N11236,N11239,N11242,N11243,N11244,N11245,N11246,N11250,N11252,N11257,
     N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,
     N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,
     N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,
     N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,
     N11316,N11317,N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,
     N11336,N11337,N11338,N11339,N11341;

  buf BUFF1_1 (N387, N1);
  buf BUFF1_2 (N388, N1);
  not NOT1_3 (N467, N57);
  and AND2_4 (N469, N134, N133);
  buf BUFF1_5 (N478, N248);
  buf BUFF1_6 (N482, N254);
  buf BUFF1_7 (N484, N257);
  buf BUFF1_8 (N486, N260);
  buf BUFF1_9 (N489, N263);
  buf BUFF1_10 (N492, N267);
  and AND4_11 (N494, N162, N172, N188, N199);
  buf BUFF1_12 (N501, N274);
  buf BUFF1_13 (N505, N280);
  buf BUFF1_14 (N507, N283);
  buf BUFF1_15 (N509, N286);
  buf BUFF1_16 (N511, N289);
  buf BUFF1_17 (N513, N293);
  buf BUFF1_18 (N515, N296);
  buf BUFF1_19 (N517, N299);
  buf BUFF1_20 (N519, N303);
  and AND4_21 (N528, N150, N184, N228, N240);
  buf BUFF1_22 (N535, N307);
  buf BUFF1_23 (N537, N310);
  buf BUFF1_24 (N539, N313);
  buf BUFF1_25 (N541, N316);
  buf BUFF1_26 (N543, N319);
  buf BUFF1_27 (N545, N322);
  buf BUFF1_28 (N547, N325);
  buf BUFF1_29 (N549, N328);
  buf BUFF1_30 (N551, N331);
  buf BUFF1_31 (N553, N334);
  buf BUFF1_32 (N556, N337);
  buf BUFF1_33 (N559, N343);
  buf BUFF1_34 (N561, N346);
  buf BUFF1_35 (N563, N349);
  buf BUFF1_36 (N565, N352);
  buf BUFF1_37 (N567, N355);
  buf BUFF1_38 (N569, N358);
  buf BUFF1_39 (N571, N361);
  buf BUFF1_40 (N573, N364);
  and AND4_41 (N575, N183, N182, N185, N186);
  and AND4_42 (N578, N210, N152, N218, N230);
  not NOT1_43 (N582, N15);
  not NOT1_44 (N585, N5);
  buf BUFF1_45 (N590, N1);
  not NOT1_46 (N593, N5);
  not NOT1_47 (N596, N5);
  not NOT1_48 (N599, N289);
  not NOT1_49 (N604, N299);
  not NOT1_50 (N609, N303);
  buf BUFF1_51 (N614, N38);
  buf BUFF1_52 (N625, N15);
  nand NAND2_53 (N628, N12, N9);
  nand NAND2_54 (N632, N12, N9);
  buf BUFF1_55 (N636, N38);
  not NOT1_56 (N641, N245);
  not NOT1_57 (N642, N248);
  buf BUFF1_58 (N643, N251);
  not NOT1_59 (N644, N251);
  not NOT1_60 (N651, N254);
  buf BUFF1_61 (N657, N106);
  not NOT1_62 (N660, N257);
  not NOT1_63 (N666, N260);
  not NOT1_64 (N672, N263);
  not NOT1_65 (N673, N267);
  not NOT1_66 (N674, N106);
  buf BUFF1_67 (N676, N18);
  buf BUFF1_68 (N682, N18);
  and AND2_69 (N688, N382, N263);
  buf BUFF1_70 (N689, N18);
  not NOT1_71 (N695, N18);
  nand NAND2_72 (N700, N382, N267);
  not NOT1_73 (N705, N271);
  not NOT1_74 (N706, N274);
  buf BUFF1_75 (N707, N277);
  not NOT1_76 (N708, N277);
  not NOT1_77 (N715, N280);
  not NOT1_78 (N721, N283);
  not NOT1_79 (N727, N286);
  not NOT1_80 (N733, N289);
  not NOT1_81 (N734, N293);
  not NOT1_82 (N742, N296);
  not NOT1_83 (N748, N299);
  not NOT1_84 (N749, N303);
  buf BUFF1_85 (N750, N367);
  not NOT1_86 (N758, N307);
  not NOT1_87 (N759, N310);
  not NOT1_88 (N762, N313);
  not NOT1_89 (N768, N316);
  not NOT1_90 (N774, N319);
  not NOT1_91 (N780, N322);
  not NOT1_92 (N786, N325);
  not NOT1_93 (N794, N328);
  not NOT1_94 (N800, N331);
  not NOT1_95 (N806, N334);
  not NOT1_96 (N812, N337);
  buf BUFF1_97 (N813, N340);
  not NOT1_98 (N814, N340);
  not NOT1_99 (N821, N343);
  not NOT1_100 (N827, N346);
  not NOT1_101 (N833, N349);
  not NOT1_102 (N839, N352);
  not NOT1_103 (N845, N355);
  not NOT1_104 (N853, N358);
  not NOT1_105 (N859, N361);
  not NOT1_106 (N865, N364);
  buf BUFF1_107 (N871, N367);
  nand NAND2_108 (N881, N467, N585);
  not NOT1_109 (N882, N528);
  not NOT1_110 (N883, N578);
  not NOT1_111 (N884, N575);
  not NOT1_112 (N885, N494);
  and AND2_113 (N886, N528, N578);
  and AND2_114 (N887, N575, N494);
  buf BUFF1_115 (N889, N590);
  buf BUFF1_116 (N945, N657);
  not NOT1_117 (N957, N688);
  and AND2_118 (N1028, N382, N641);
  nand NAND2_119 (N1029, N382, N705);
  and AND2_120 (N1109, N469, N596);
  nand NAND2_121 (N1110, N242, N593);
  not NOT1_122 (N1111, N625);
  nand NAND2_123 (N1112, N242, N593);
  nand NAND2_124 (N1113, N469, N596);
  not NOT1_125 (N1114, N625);
  not NOT1_126 (N1115, N871);
  buf BUFF1_127 (N1116, N590);
  buf BUFF1_128 (N1119, N628);
  buf BUFF1_129 (N1125, N682);
  buf BUFF1_130 (N1132, N628);
  buf BUFF1_131 (N1136, N682);
  buf BUFF1_132 (N1141, N628);
  buf BUFF1_133 (N1147, N682);
  buf BUFF1_134 (N1154, N632);
  buf BUFF1_135 (N1160, N676);
  and AND2_136 (N1167, N700, N614);
  and AND2_137 (N1174, N700, N614);
  buf BUFF1_138 (N1175, N682);
  buf BUFF1_139 (N1182, N676);
  not NOT1_140 (N1189, N657);
  not NOT1_141 (N1194, N676);
  not NOT1_142 (N1199, N682);
  not NOT1_143 (N1206, N689);
  buf BUFF1_144 (N1211, N695);
  not NOT1_145 (N1218, N750);
  not NOT1_146 (N1222, N1028);
  buf BUFF1_147 (N1227, N632);
  buf BUFF1_148 (N1233, N676);
  buf BUFF1_149 (N1240, N632);
  buf BUFF1_150 (N1244, N676);
  buf BUFF1_151 (N1249, N689);
  buf BUFF1_152 (N1256, N689);
  buf BUFF1_153 (N1263, N695);
  buf BUFF1_154 (N1270, N689);
  buf BUFF1_155 (N1277, N689);
  buf BUFF1_156 (N1284, N700);
  buf BUFF1_157 (N1287, N614);
  buf BUFF1_158 (N1290, N666);
  buf BUFF1_159 (N1293, N660);
  buf BUFF1_160 (N1296, N651);
  buf BUFF1_161 (N1299, N614);
  buf BUFF1_162 (N1302, N644);
  buf BUFF1_163 (N1305, N700);
  buf BUFF1_164 (N1308, N614);
  buf BUFF1_165 (N1311, N614);
  buf BUFF1_166 (N1314, N666);
  buf BUFF1_167 (N1317, N660);
  buf BUFF1_168 (N1320, N651);
  buf BUFF1_169 (N1323, N644);
  buf BUFF1_170 (N1326, N609);
  buf BUFF1_171 (N1329, N604);
  buf BUFF1_172 (N1332, N742);
  buf BUFF1_173 (N1335, N599);
  buf BUFF1_174 (N1338, N727);
  buf BUFF1_175 (N1341, N721);
  buf BUFF1_176 (N1344, N715);
  buf BUFF1_177 (N1347, N734);
  buf BUFF1_178 (N1350, N708);
  buf BUFF1_179 (N1353, N609);
  buf BUFF1_180 (N1356, N604);
  buf BUFF1_181 (N1359, N742);
  buf BUFF1_182 (N1362, N734);
  buf BUFF1_183 (N1365, N599);
  buf BUFF1_184 (N1368, N727);
  buf BUFF1_185 (N1371, N721);
  buf BUFF1_186 (N1374, N715);
  buf BUFF1_187 (N1377, N708);
  buf BUFF1_188 (N1380, N806);
  buf BUFF1_189 (N1383, N800);
  buf BUFF1_190 (N1386, N794);
  buf BUFF1_191 (N1389, N786);
  buf BUFF1_192 (N1392, N780);
  buf BUFF1_193 (N1395, N774);
  buf BUFF1_194 (N1398, N768);
  buf BUFF1_195 (N1401, N762);
  buf BUFF1_196 (N1404, N806);
  buf BUFF1_197 (N1407, N800);
  buf BUFF1_198 (N1410, N794);
  buf BUFF1_199 (N1413, N780);
  buf BUFF1_200 (N1416, N774);
  buf BUFF1_201 (N1419, N768);
  buf BUFF1_202 (N1422, N762);
  buf BUFF1_203 (N1425, N786);
  buf BUFF1_204 (N1428, N636);
  buf BUFF1_205 (N1431, N636);
  buf BUFF1_206 (N1434, N865);
  buf BUFF1_207 (N1437, N859);
  buf BUFF1_208 (N1440, N853);
  buf BUFF1_209 (N1443, N845);
  buf BUFF1_210 (N1446, N839);
  buf BUFF1_211 (N1449, N833);
  buf BUFF1_212 (N1452, N827);
  buf BUFF1_213 (N1455, N821);
  buf BUFF1_214 (N1458, N814);
  buf BUFF1_215 (N1461, N865);
  buf BUFF1_216 (N1464, N859);
  buf BUFF1_217 (N1467, N853);
  buf BUFF1_218 (N1470, N839);
  buf BUFF1_219 (N1473, N833);
  buf BUFF1_220 (N1476, N827);
  buf BUFF1_221 (N1479, N821);
  buf BUFF1_222 (N1482, N845);
  buf BUFF1_223 (N1485, N814);
  not NOT1_224 (N1489, N1109);
  buf BUFF1_225 (N1490, N1116);
  and AND2_226 (N1537, N957, N614);
  and AND2_227 (N1551, N614, N957);
  and AND2_228 (N1649, N1029, N636);
  buf BUFF1_229 (N1703, N957);
  nor NOR2_230 (N1708, N957, N614);
  buf BUFF1_231 (N1713, N957);
  nor NOR2_232 (N1721, N614, N957);
  buf BUFF1_233 (N1758, N1029);
  and AND2_234 (N1781, N163, N1116);
  and AND2_235 (N1782, N170, N1125);
  not NOT1_236 (N1783, N1125);
  not NOT1_237 (N1789, N1136);
  and AND2_238 (N1793, N169, N1125);
  and AND2_239 (N1794, N168, N1125);
  and AND2_240 (N1795, N167, N1125);
  and AND2_241 (N1796, N166, N1136);
  and AND2_242 (N1797, N165, N1136);
  and AND2_243 (N1798, N164, N1136);
  not NOT1_244 (N1799, N1147);
  not NOT1_245 (N1805, N1160);
  and AND2_246 (N1811, N177, N1147);
  and AND2_247 (N1812, N176, N1147);
  and AND2_248 (N1813, N175, N1147);
  and AND2_249 (N1814, N174, N1147);
  and AND2_250 (N1815, N173, N1147);
  and AND2_251 (N1816, N157, N1160);
  and AND2_252 (N1817, N156, N1160);
  and AND2_253 (N1818, N155, N1160);
  and AND2_254 (N1819, N154, N1160);
  and AND2_255 (N1820, N153, N1160);
  not NOT1_256 (N1821, N1284);
  not NOT1_257 (N1822, N1287);
  not NOT1_258 (N1828, N1290);
  not NOT1_259 (N1829, N1293);
  not NOT1_260 (N1830, N1296);
  not NOT1_261 (N1832, N1299);
  not NOT1_262 (N1833, N1302);
  not NOT1_263 (N1834, N1305);
  not NOT1_264 (N1835, N1308);
  not NOT1_265 (N1839, N1311);
  not NOT1_266 (N1840, N1314);
  not NOT1_267 (N1841, N1317);
  not NOT1_268 (N1842, N1320);
  not NOT1_269 (N1843, N1323);
  not NOT1_270 (N1845, N1175);
  not NOT1_271 (N1851, N1182);
  and AND2_272 (N1857, N181, N1175);
  and AND2_273 (N1858, N171, N1175);
  and AND2_274 (N1859, N180, N1175);
  and AND2_275 (N1860, N179, N1175);
  and AND2_276 (N1861, N178, N1175);
  and AND2_277 (N1862, N161, N1182);
  and AND2_278 (N1863, N151, N1182);
  and AND2_279 (N1864, N160, N1182);
  and AND2_280 (N1865, N159, N1182);
  and AND2_281 (N1866, N158, N1182);
  not NOT1_282 (N1867, N1326);
  not NOT1_283 (N1868, N1329);
  not NOT1_284 (N1869, N1332);
  not NOT1_285 (N1870, N1335);
  not NOT1_286 (N1871, N1338);
  not NOT1_287 (N1872, N1341);
  not NOT1_288 (N1873, N1344);
  not NOT1_289 (N1874, N1347);
  not NOT1_290 (N1875, N1350);
  not NOT1_291 (N1876, N1353);
  not NOT1_292 (N1877, N1356);
  not NOT1_293 (N1878, N1359);
  not NOT1_294 (N1879, N1362);
  not NOT1_295 (N1880, N1365);
  not NOT1_296 (N1881, N1368);
  not NOT1_297 (N1882, N1371);
  not NOT1_298 (N1883, N1374);
  not NOT1_299 (N1884, N1377);
  buf BUFF1_300 (N1885, N1199);
  buf BUFF1_301 (N1892, N1194);
  buf BUFF1_302 (N1899, N1199);
  buf BUFF1_303 (N1906, N1194);
  not NOT1_304 (N1913, N1211);
  buf BUFF1_305 (N1919, N1194);
  and AND2_306 (N1926, N44, N1211);
  and AND2_307 (N1927, N41, N1211);
  and AND2_308 (N1928, N29, N1211);
  and AND2_309 (N1929, N26, N1211);
  and AND2_310 (N1930, N23, N1211);
  not NOT1_311 (N1931, N1380);
  not NOT1_312 (N1932, N1383);
  not NOT1_313 (N1933, N1386);
  not NOT1_314 (N1934, N1389);
  not NOT1_315 (N1935, N1392);
  not NOT1_316 (N1936, N1395);
  not NOT1_317 (N1937, N1398);
  not NOT1_318 (N1938, N1401);
  not NOT1_319 (N1939, N1404);
  not NOT1_320 (N1940, N1407);
  not NOT1_321 (N1941, N1410);
  not NOT1_322 (N1942, N1413);
  not NOT1_323 (N1943, N1416);
  not NOT1_324 (N1944, N1419);
  not NOT1_325 (N1945, N1422);
  not NOT1_326 (N1946, N1425);
  not NOT1_327 (N1947, N1233);
  not NOT1_328 (N1953, N1244);
  and AND2_329 (N1957, N209, N1233);
  and AND2_330 (N1958, N216, N1233);
  and AND2_331 (N1959, N215, N1233);
  and AND2_332 (N1960, N214, N1233);
  and AND2_333 (N1961, N213, N1244);
  and AND2_334 (N1962, N212, N1244);
  and AND2_335 (N1963, N211, N1244);
  not NOT1_336 (N1965, N1428);
  and AND2_337 (N1966, N1222, N636);
  not NOT1_338 (N1967, N1431);
  not NOT1_339 (N1968, N1434);
  not NOT1_340 (N1969, N1437);
  not NOT1_341 (N1970, N1440);
  not NOT1_342 (N1971, N1443);
  not NOT1_343 (N1972, N1446);
  not NOT1_344 (N1973, N1449);
  not NOT1_345 (N1974, N1452);
  not NOT1_346 (N1975, N1455);
  not NOT1_347 (N1976, N1458);
  not NOT1_348 (N1977, N1249);
  not NOT1_349 (N1983, N1256);
  and AND2_350 (N1989, N642, N1249);
  and AND2_351 (N1990, N644, N1249);
  and AND2_352 (N1991, N651, N1249);
  and AND2_353 (N1992, N674, N1249);
  and AND2_354 (N1993, N660, N1249);
  and AND2_355 (N1994, N666, N1256);
  and AND2_356 (N1995, N672, N1256);
  and AND2_357 (N1996, N673, N1256);
  not NOT1_358 (N1997, N1263);
  buf BUFF1_359 (N2003, N1194);
  and AND2_360 (N2010, N47, N1263);
  and AND2_361 (N2011, N35, N1263);
  and AND2_362 (N2012, N32, N1263);
  and AND2_363 (N2013, N50, N1263);
  and AND2_364 (N2014, N66, N1263);
  not NOT1_365 (N2015, N1461);
  not NOT1_366 (N2016, N1464);
  not NOT1_367 (N2017, N1467);
  not NOT1_368 (N2018, N1470);
  not NOT1_369 (N2019, N1473);
  not NOT1_370 (N2020, N1476);
  not NOT1_371 (N2021, N1479);
  not NOT1_372 (N2022, N1482);
  not NOT1_373 (N2023, N1485);
  buf BUFF1_374 (N2024, N1206);
  buf BUFF1_375 (N2031, N1206);
  buf BUFF1_376 (N2038, N1206);
  buf BUFF1_377 (N2045, N1206);
  not NOT1_378 (N2052, N1270);
  not NOT1_379 (N2058, N1277);
  and AND2_380 (N2064, N706, N1270);
  and AND2_381 (N2065, N708, N1270);
  and AND2_382 (N2066, N715, N1270);
  and AND2_383 (N2067, N721, N1270);
  and AND2_384 (N2068, N727, N1270);
  and AND2_385 (N2069, N733, N1277);
  and AND2_386 (N2070, N734, N1277);
  and AND2_387 (N2071, N742, N1277);
  and AND2_388 (N2072, N748, N1277);
  and AND2_389 (N2073, N749, N1277);
  buf BUFF1_390 (N2074, N1189);
  buf BUFF1_391 (N2081, N1189);
  buf BUFF1_392 (N2086, N1222);
  nand NAND2_393 (N2107, N1287, N1821);
  nand NAND2_394 (N2108, N1284, N1822);
  not NOT1_395 (N2110, N1703);
  nand NAND2_396 (N2111, N1703, N1832);
  nand NAND2_397 (N2112, N1308, N1834);
  nand NAND2_398 (N2113, N1305, N1835);
  not NOT1_399 (N2114, N1713);
  nand NAND2_400 (N2115, N1713, N1839);
  not NOT1_401 (N2117, N1721);
  not NOT1_402 (N2171, N1758);
  nand NAND2_403 (N2172, N1758, N1965);
  not NOT1_404 (N2230, N1708);
  buf BUFF1_405 (N2231, N1537);
  buf BUFF1_406 (N2235, N1551);
  or OR2_407 (N2239, N1783, N1782);
  or OR2_408 (N2240, N1783, N1125);
  or OR2_409 (N2241, N1783, N1793);
  or OR2_410 (N2242, N1783, N1794);
  or OR2_411 (N2243, N1783, N1795);
  or OR2_412 (N2244, N1789, N1796);
  or OR2_413 (N2245, N1789, N1797);
  or OR2_414 (N2246, N1789, N1798);
  or OR2_415 (N2247, N1799, N1811);
  or OR2_416 (N2248, N1799, N1812);
  or OR2_417 (N2249, N1799, N1813);
  or OR2_418 (N2250, N1799, N1814);
  or OR2_419 (N2251, N1799, N1815);
  or OR2_420 (N2252, N1805, N1816);
  or OR2_421 (N2253, N1805, N1817);
  or OR2_422 (N2254, N1805, N1818);
  or OR2_423 (N2255, N1805, N1819);
  or OR2_424 (N2256, N1805, N1820);
  nand NAND2_425 (N2257, N2107, N2108);
  not NOT1_426 (N2267, N2074);
  nand NAND2_427 (N2268, N1299, N2110);
  nand NAND2_428 (N2269, N2112, N2113);
  nand NAND2_429 (N2274, N1311, N2114);
  not NOT1_430 (N2275, N2081);
  and AND2_431 (N2277, N141, N1845);
  and AND2_432 (N2278, N147, N1845);
  and AND2_433 (N2279, N138, N1845);
  and AND2_434 (N2280, N144, N1845);
  and AND2_435 (N2281, N135, N1845);
  and AND2_436 (N2282, N141, N1851);
  and AND2_437 (N2283, N147, N1851);
  and AND2_438 (N2284, N138, N1851);
  and AND2_439 (N2285, N144, N1851);
  and AND2_440 (N2286, N135, N1851);
  not NOT1_441 (N2287, N1885);
  not NOT1_442 (N2293, N1892);
  and AND2_443 (N2299, N103, N1885);
  and AND2_444 (N2300, N130, N1885);
  and AND2_445 (N2301, N127, N1885);
  and AND2_446 (N2302, N124, N1885);
  and AND2_447 (N2303, N100, N1885);
  and AND2_448 (N2304, N103, N1892);
  and AND2_449 (N2305, N130, N1892);
  and AND2_450 (N2306, N127, N1892);
  and AND2_451 (N2307, N124, N1892);
  and AND2_452 (N2308, N100, N1892);
  not NOT1_453 (N2309, N1899);
  not NOT1_454 (N2315, N1906);
  and AND2_455 (N2321, N115, N1899);
  and AND2_456 (N2322, N118, N1899);
  and AND2_457 (N2323, N97, N1899);
  and AND2_458 (N2324, N94, N1899);
  and AND2_459 (N2325, N121, N1899);
  and AND2_460 (N2326, N115, N1906);
  and AND2_461 (N2327, N118, N1906);
  and AND2_462 (N2328, N97, N1906);
  and AND2_463 (N2329, N94, N1906);
  and AND2_464 (N2330, N121, N1906);
  not NOT1_465 (N2331, N1919);
  and AND2_466 (N2337, N208, N1913);
  and AND2_467 (N2338, N198, N1913);
  and AND2_468 (N2339, N207, N1913);
  and AND2_469 (N2340, N206, N1913);
  and AND2_470 (N2341, N205, N1913);
  and AND2_471 (N2342, N44, N1919);
  and AND2_472 (N2343, N41, N1919);
  and AND2_473 (N2344, N29, N1919);
  and AND2_474 (N2345, N26, N1919);
  and AND2_475 (N2346, N23, N1919);
  or OR2_476 (N2347, N1947, N1233);
  or OR2_477 (N2348, N1947, N1957);
  or OR2_478 (N2349, N1947, N1958);
  or OR2_479 (N2350, N1947, N1959);
  or OR2_480 (N2351, N1947, N1960);
  or OR2_481 (N2352, N1953, N1961);
  or OR2_482 (N2353, N1953, N1962);
  or OR2_483 (N2354, N1953, N1963);
  nand NAND2_484 (N2355, N1428, N2171);
  not NOT1_485 (N2356, N2086);
  nand NAND2_486 (N2357, N2086, N1967);
  and AND2_487 (N2358, N114, N1977);
  and AND2_488 (N2359, N113, N1977);
  and AND2_489 (N2360, N111, N1977);
  and AND2_490 (N2361, N87, N1977);
  and AND2_491 (N2362, N112, N1977);
  and AND2_492 (N2363, N88, N1983);
  and AND2_493 (N2364, N245, N1983);
  and AND2_494 (N2365, N271, N1983);
  and AND2_495 (N2366, N759, N1983);
  and AND2_496 (N2367, N70, N1983);
  not NOT1_497 (N2368, N2003);
  and AND2_498 (N2374, N193, N1997);
  and AND2_499 (N2375, N192, N1997);
  and AND2_500 (N2376, N191, N1997);
  and AND2_501 (N2377, N190, N1997);
  and AND2_502 (N2378, N189, N1997);
  and AND2_503 (N2379, N47, N2003);
  and AND2_504 (N2380, N35, N2003);
  and AND2_505 (N2381, N32, N2003);
  and AND2_506 (N2382, N50, N2003);
  and AND2_507 (N2383, N66, N2003);
  not NOT1_508 (N2384, N2024);
  not NOT1_509 (N2390, N2031);
  and AND2_510 (N2396, N58, N2024);
  and AND2_511 (N2397, N77, N2024);
  and AND2_512 (N2398, N78, N2024);
  and AND2_513 (N2399, N59, N2024);
  and AND2_514 (N2400, N81, N2024);
  and AND2_515 (N2401, N80, N2031);
  and AND2_516 (N2402, N79, N2031);
  and AND2_517 (N2403, N60, N2031);
  and AND2_518 (N2404, N61, N2031);
  and AND2_519 (N2405, N62, N2031);
  not NOT1_520 (N2406, N2038);
  not NOT1_521 (N2412, N2045);
  and AND2_522 (N2418, N69, N2038);
  and AND2_523 (N2419, N70, N2038);
  and AND2_524 (N2420, N74, N2038);
  and AND2_525 (N2421, N76, N2038);
  and AND2_526 (N2422, N75, N2038);
  and AND2_527 (N2423, N73, N2045);
  and AND2_528 (N2424, N53, N2045);
  and AND2_529 (N2425, N54, N2045);
  and AND2_530 (N2426, N55, N2045);
  and AND2_531 (N2427, N56, N2045);
  and AND2_532 (N2428, N82, N2052);
  and AND2_533 (N2429, N65, N2052);
  and AND2_534 (N2430, N83, N2052);
  and AND2_535 (N2431, N84, N2052);
  and AND2_536 (N2432, N85, N2052);
  and AND2_537 (N2433, N64, N2058);
  and AND2_538 (N2434, N63, N2058);
  and AND2_539 (N2435, N86, N2058);
  and AND2_540 (N2436, N109, N2058);
  and AND2_541 (N2437, N110, N2058);
  and AND2_542 (N2441, N2239, N1119);
  and AND2_543 (N2442, N2240, N1119);
  and AND2_544 (N2446, N2241, N1119);
  and AND2_545 (N2450, N2242, N1119);
  and AND2_546 (N2454, N2243, N1119);
  and AND2_547 (N2458, N2244, N1132);
  and AND2_548 (N2462, N2247, N1141);
  and AND2_549 (N2466, N2248, N1141);
  and AND2_550 (N2470, N2249, N1141);
  and AND2_551 (N2474, N2250, N1141);
  and AND2_552 (N2478, N2251, N1141);
  and AND2_553 (N2482, N2252, N1154);
  and AND2_554 (N2488, N2253, N1154);
  and AND2_555 (N2496, N2254, N1154);
  and AND2_556 (N2502, N2255, N1154);
  and AND2_557 (N2508, N2256, N1154);
  nand NAND2_558 (N2523, N2268, N2111);
  nand NAND2_559 (N2533, N2274, N2115);
  not NOT1_560 (N2537, N2235);
  or OR2_561 (N2538, N2278, N1858);
  or OR2_562 (N2542, N2279, N1859);
  or OR2_563 (N2546, N2280, N1860);
  or OR2_564 (N2550, N2281, N1861);
  or OR2_565 (N2554, N2283, N1863);
  or OR2_566 (N2561, N2284, N1864);
  or OR2_567 (N2567, N2285, N1865);
  or OR2_568 (N2573, N2286, N1866);
  or OR2_569 (N2604, N2338, N1927);
  or OR2_570 (N2607, N2339, N1928);
  or OR2_571 (N2611, N2340, N1929);
  or OR2_572 (N2615, N2341, N1930);
  and AND2_573 (N2619, N2348, N1227);
  and AND2_574 (N2626, N2349, N1227);
  and AND2_575 (N2632, N2350, N1227);
  and AND2_576 (N2638, N2351, N1227);
  and AND2_577 (N2644, N2352, N1240);
  nand NAND2_578 (N2650, N2355, N2172);
  nand NAND2_579 (N2653, N1431, N2356);
  or OR2_580 (N2654, N2359, N1990);
  or OR2_581 (N2658, N2360, N1991);
  or OR2_582 (N2662, N2361, N1992);
  or OR2_583 (N2666, N2362, N1993);
  or OR2_584 (N2670, N2363, N1994);
  or OR2_585 (N2674, N2366, N1256);
  or OR2_586 (N2680, N2367, N1256);
  or OR2_587 (N2688, N2374, N2010);
  or OR2_588 (N2692, N2375, N2011);
  or OR2_589 (N2696, N2376, N2012);
  or OR2_590 (N2700, N2377, N2013);
  or OR2_591 (N2704, N2378, N2014);
  and AND2_592 (N2728, N2347, N1227);
  or OR2_593 (N2729, N2429, N2065);
  or OR2_594 (N2733, N2430, N2066);
  or OR2_595 (N2737, N2431, N2067);
  or OR2_596 (N2741, N2432, N2068);
  or OR2_597 (N2745, N2433, N2069);
  or OR2_598 (N2749, N2434, N2070);
  or OR2_599 (N2753, N2435, N2071);
  or OR2_600 (N2757, N2436, N2072);
  or OR2_601 (N2761, N2437, N2073);
  not NOT1_602 (N2765, N2231);
  and AND2_603 (N2766, N2354, N1240);
  and AND2_604 (N2769, N2353, N1240);
  and AND2_605 (N2772, N2246, N1132);
  and AND2_606 (N2775, N2245, N1132);
  or OR2_607 (N2778, N2282, N1862);
  or OR2_608 (N2781, N2358, N1989);
  or OR2_609 (N2784, N2365, N1996);
  or OR2_610 (N2787, N2364, N1995);
  or OR2_611 (N2790, N2337, N1926);
  or OR2_612 (N2793, N2277, N1857);
  or OR2_613 (N2796, N2428, N2064);
  and AND2_614 (N2866, N2257, N1537);
  and AND2_615 (N2867, N2257, N1537);
  and AND2_616 (N2868, N2257, N1537);
  and AND2_617 (N2869, N2257, N1537);
  and AND2_618 (N2878, N2269, N1551);
  and AND2_619 (N2913, N204, N2287);
  and AND2_620 (N2914, N203, N2287);
  and AND2_621 (N2915, N202, N2287);
  and AND2_622 (N2916, N201, N2287);
  and AND2_623 (N2917, N200, N2287);
  and AND2_624 (N2918, N235, N2293);
  and AND2_625 (N2919, N234, N2293);
  and AND2_626 (N2920, N233, N2293);
  and AND2_627 (N2921, N232, N2293);
  and AND2_628 (N2922, N231, N2293);
  and AND2_629 (N2923, N197, N2309);
  and AND2_630 (N2924, N187, N2309);
  and AND2_631 (N2925, N196, N2309);
  and AND2_632 (N2926, N195, N2309);
  and AND2_633 (N2927, N194, N2309);
  and AND2_634 (N2928, N227, N2315);
  and AND2_635 (N2929, N217, N2315);
  and AND2_636 (N2930, N226, N2315);
  and AND2_637 (N2931, N225, N2315);
  and AND2_638 (N2932, N224, N2315);
  and AND2_639 (N2933, N239, N2331);
  and AND2_640 (N2934, N229, N2331);
  and AND2_641 (N2935, N238, N2331);
  and AND2_642 (N2936, N237, N2331);
  and AND2_643 (N2937, N236, N2331);
  nand NAND2_644 (N2988, N2653, N2357);
  and AND2_645 (N3005, N223, N2368);
  and AND2_646 (N3006, N222, N2368);
  and AND2_647 (N3007, N221, N2368);
  and AND2_648 (N3008, N220, N2368);
  and AND2_649 (N3009, N219, N2368);
  and AND2_650 (N3020, N812, N2384);
  and AND2_651 (N3021, N814, N2384);
  and AND2_652 (N3022, N821, N2384);
  and AND2_653 (N3023, N827, N2384);
  and AND2_654 (N3024, N833, N2384);
  and AND2_655 (N3025, N839, N2390);
  and AND2_656 (N3026, N845, N2390);
  and AND2_657 (N3027, N853, N2390);
  and AND2_658 (N3028, N859, N2390);
  and AND2_659 (N3029, N865, N2390);
  and AND2_660 (N3032, N758, N2406);
  and AND2_661 (N3033, N759, N2406);
  and AND2_662 (N3034, N762, N2406);
  and AND2_663 (N3035, N768, N2406);
  and AND2_664 (N3036, N774, N2406);
  and AND2_665 (N3037, N780, N2412);
  and AND2_666 (N3038, N786, N2412);
  and AND2_667 (N3039, N794, N2412);
  and AND2_668 (N3040, N800, N2412);
  and AND2_669 (N3041, N806, N2412);
  buf BUFF1_670 (N3061, N2257);
  buf BUFF1_671 (N3064, N2257);
  buf BUFF1_672 (N3067, N2269);
  buf BUFF1_673 (N3070, N2269);
  not NOT1_674 (N3073, N2728);
  not NOT1_675 (N3080, N2441);
  and AND2_676 (N3096, N666, N2644);
  and AND2_677 (N3097, N660, N2638);
  and AND2_678 (N3101, N1189, N2632);
  and AND2_679 (N3107, N651, N2626);
  and AND2_680 (N3114, N644, N2619);
  and AND2_681 (N3122, N2523, N2257);
  or OR2_682 (N3126, N1167, N2866);
  and AND2_683 (N3130, N2523, N2257);
  or OR2_684 (N3131, N1167, N2869);
  and AND2_685 (N3134, N2523, N2257);
  not NOT1_686 (N3135, N2533);
  and AND2_687 (N3136, N666, N2644);
  and AND2_688 (N3137, N660, N2638);
  and AND2_689 (N3140, N1189, N2632);
  and AND2_690 (N3144, N651, N2626);
  and AND2_691 (N3149, N644, N2619);
  and AND2_692 (N3155, N2533, N2269);
  or OR2_693 (N3159, N1174, N2878);
  not NOT1_694 (N3167, N2778);
  and AND2_695 (N3168, N609, N2508);
  and AND2_696 (N3169, N604, N2502);
  and AND2_697 (N3173, N742, N2496);
  and AND2_698 (N3178, N734, N2488);
  and AND2_699 (N3184, N599, N2482);
  and AND2_700 (N3185, N727, N2573);
  and AND2_701 (N3189, N721, N2567);
  and AND2_702 (N3195, N715, N2561);
  and AND2_703 (N3202, N708, N2554);
  and AND2_704 (N3210, N609, N2508);
  and AND2_705 (N3211, N604, N2502);
  and AND2_706 (N3215, N742, N2496);
  and AND2_707 (N3221, N2488, N734);
  and AND2_708 (N3228, N599, N2482);
  and AND2_709 (N3229, N727, N2573);
  and AND2_710 (N3232, N721, N2567);
  and AND2_711 (N3236, N715, N2561);
  and AND2_712 (N3241, N708, N2554);
  or OR2_713 (N3247, N2913, N2299);
  or OR2_714 (N3251, N2914, N2300);
  or OR2_715 (N3255, N2915, N2301);
  or OR2_716 (N3259, N2916, N2302);
  or OR2_717 (N3263, N2917, N2303);
  or OR2_718 (N3267, N2918, N2304);
  or OR2_719 (N3273, N2919, N2305);
  or OR2_720 (N3281, N2920, N2306);
  or OR2_721 (N3287, N2921, N2307);
  or OR2_722 (N3293, N2922, N2308);
  or OR2_723 (N3299, N2924, N2322);
  or OR2_724 (N3303, N2925, N2323);
  or OR2_725 (N3307, N2926, N2324);
  or OR2_726 (N3311, N2927, N2325);
  or OR2_727 (N3315, N2929, N2327);
  or OR2_728 (N3322, N2930, N2328);
  or OR2_729 (N3328, N2931, N2329);
  or OR2_730 (N3334, N2932, N2330);
  or OR2_731 (N3340, N2934, N2343);
  or OR2_732 (N3343, N2935, N2344);
  or OR2_733 (N3349, N2936, N2345);
  or OR2_734 (N3355, N2937, N2346);
  and AND2_735 (N3361, N2761, N2478);
  and AND2_736 (N3362, N2757, N2474);
  and AND2_737 (N3363, N2753, N2470);
  and AND2_738 (N3364, N2749, N2466);
  and AND2_739 (N3365, N2745, N2462);
  and AND2_740 (N3366, N2741, N2550);
  and AND2_741 (N3367, N2737, N2546);
  and AND2_742 (N3368, N2733, N2542);
  and AND2_743 (N3369, N2729, N2538);
  and AND2_744 (N3370, N2670, N2458);
  and AND2_745 (N3371, N2666, N2454);
  and AND2_746 (N3372, N2662, N2450);
  and AND2_747 (N3373, N2658, N2446);
  and AND2_748 (N3374, N2654, N2442);
  and AND2_749 (N3375, N2988, N2650);
  and AND2_750 (N3379, N2650, N1966);
  not NOT1_751 (N3380, N2781);
  and AND2_752 (N3381, N695, N2604);
  or OR2_753 (N3384, N3005, N2379);
  or OR2_754 (N3390, N3006, N2380);
  or OR2_755 (N3398, N3007, N2381);
  or OR2_756 (N3404, N3008, N2382);
  or OR2_757 (N3410, N3009, N2383);
  or OR2_758 (N3416, N3021, N2397);
  or OR2_759 (N3420, N3022, N2398);
  or OR2_760 (N3424, N3023, N2399);
  or OR2_761 (N3428, N3024, N2400);
  or OR2_762 (N3432, N3025, N2401);
  or OR2_763 (N3436, N3026, N2402);
  or OR2_764 (N3440, N3027, N2403);
  or OR2_765 (N3444, N3028, N2404);
  or OR2_766 (N3448, N3029, N2405);
  not NOT1_767 (N3452, N2790);
  not NOT1_768 (N3453, N2793);
  or OR2_769 (N3454, N3034, N2420);
  or OR2_770 (N3458, N3035, N2421);
  or OR2_771 (N3462, N3036, N2422);
  or OR2_772 (N3466, N3037, N2423);
  or OR2_773 (N3470, N3038, N2424);
  or OR2_774 (N3474, N3039, N2425);
  or OR2_775 (N3478, N3040, N2426);
  or OR2_776 (N3482, N3041, N2427);
  not NOT1_777 (N3486, N2796);
  buf BUFF1_778 (N3487, N2644);
  buf BUFF1_779 (N3490, N2638);
  buf BUFF1_780 (N3493, N2632);
  buf BUFF1_781 (N3496, N2626);
  buf BUFF1_782 (N3499, N2619);
  buf BUFF1_783 (N3502, N2523);
  nor NOR2_784 (N3507, N1167, N2868);
  buf BUFF1_785 (N3510, N2523);
  nor NOR2_786 (N3515, N644, N2619);
  buf BUFF1_787 (N3518, N2644);
  buf BUFF1_788 (N3521, N2638);
  buf BUFF1_789 (N3524, N2632);
  buf BUFF1_790 (N3527, N2626);
  buf BUFF1_791 (N3530, N2619);
  buf BUFF1_792 (N3535, N2619);
  buf BUFF1_793 (N3539, N2632);
  buf BUFF1_794 (N3542, N2626);
  buf BUFF1_795 (N3545, N2644);
  buf BUFF1_796 (N3548, N2638);
  not NOT1_797 (N3551, N2766);
  not NOT1_798 (N3552, N2769);
  buf BUFF1_799 (N3553, N2442);
  buf BUFF1_800 (N3557, N2450);
  buf BUFF1_801 (N3560, N2446);
  buf BUFF1_802 (N3563, N2458);
  buf BUFF1_803 (N3566, N2454);
  not NOT1_804 (N3569, N2772);
  not NOT1_805 (N3570, N2775);
  buf BUFF1_806 (N3571, N2554);
  buf BUFF1_807 (N3574, N2567);
  buf BUFF1_808 (N3577, N2561);
  buf BUFF1_809 (N3580, N2482);
  buf BUFF1_810 (N3583, N2573);
  buf BUFF1_811 (N3586, N2496);
  buf BUFF1_812 (N3589, N2488);
  buf BUFF1_813 (N3592, N2508);
  buf BUFF1_814 (N3595, N2502);
  buf BUFF1_815 (N3598, N2508);
  buf BUFF1_816 (N3601, N2502);
  buf BUFF1_817 (N3604, N2496);
  buf BUFF1_818 (N3607, N2482);
  buf BUFF1_819 (N3610, N2573);
  buf BUFF1_820 (N3613, N2567);
  buf BUFF1_821 (N3616, N2561);
  buf BUFF1_822 (N3619, N2488);
  buf BUFF1_823 (N3622, N2554);
  nor NOR2_824 (N3625, N734, N2488);
  nor NOR2_825 (N3628, N708, N2554);
  buf BUFF1_826 (N3631, N2508);
  buf BUFF1_827 (N3634, N2502);
  buf BUFF1_828 (N3637, N2496);
  buf BUFF1_829 (N3640, N2488);
  buf BUFF1_830 (N3643, N2482);
  buf BUFF1_831 (N3646, N2573);
  buf BUFF1_832 (N3649, N2567);
  buf BUFF1_833 (N3652, N2561);
  buf BUFF1_834 (N3655, N2554);
  nor NOR2_835 (N3658, N2488, N734);
  buf BUFF1_836 (N3661, N2674);
  buf BUFF1_837 (N3664, N2674);
  buf BUFF1_838 (N3667, N2761);
  buf BUFF1_839 (N3670, N2478);
  buf BUFF1_840 (N3673, N2757);
  buf BUFF1_841 (N3676, N2474);
  buf BUFF1_842 (N3679, N2753);
  buf BUFF1_843 (N3682, N2470);
  buf BUFF1_844 (N3685, N2745);
  buf BUFF1_845 (N3688, N2462);
  buf BUFF1_846 (N3691, N2741);
  buf BUFF1_847 (N3694, N2550);
  buf BUFF1_848 (N3697, N2737);
  buf BUFF1_849 (N3700, N2546);
  buf BUFF1_850 (N3703, N2733);
  buf BUFF1_851 (N3706, N2542);
  buf BUFF1_852 (N3709, N2749);
  buf BUFF1_853 (N3712, N2466);
  buf BUFF1_854 (N3715, N2729);
  buf BUFF1_855 (N3718, N2538);
  buf BUFF1_856 (N3721, N2704);
  buf BUFF1_857 (N3724, N2700);
  buf BUFF1_858 (N3727, N2696);
  buf BUFF1_859 (N3730, N2688);
  buf BUFF1_860 (N3733, N2692);
  buf BUFF1_861 (N3736, N2670);
  buf BUFF1_862 (N3739, N2458);
  buf BUFF1_863 (N3742, N2666);
  buf BUFF1_864 (N3745, N2454);
  buf BUFF1_865 (N3748, N2662);
  buf BUFF1_866 (N3751, N2450);
  buf BUFF1_867 (N3754, N2658);
  buf BUFF1_868 (N3757, N2446);
  buf BUFF1_869 (N3760, N2654);
  buf BUFF1_870 (N3763, N2442);
  buf BUFF1_871 (N3766, N2654);
  buf BUFF1_872 (N3769, N2662);
  buf BUFF1_873 (N3772, N2658);
  buf BUFF1_874 (N3775, N2670);
  buf BUFF1_875 (N3778, N2666);
  not NOT1_876 (N3781, N2784);
  not NOT1_877 (N3782, N2787);
  or OR2_878 (N3783, N2928, N2326);
  or OR2_879 (N3786, N2933, N2342);
  or OR2_880 (N3789, N2923, N2321);
  buf BUFF1_881 (N3792, N2688);
  buf BUFF1_882 (N3795, N2696);
  buf BUFF1_883 (N3798, N2692);
  buf BUFF1_884 (N3801, N2704);
  buf BUFF1_885 (N3804, N2700);
  buf BUFF1_886 (N3807, N2604);
  buf BUFF1_887 (N3810, N2611);
  buf BUFF1_888 (N3813, N2607);
  buf BUFF1_889 (N3816, N2615);
  buf BUFF1_890 (N3819, N2538);
  buf BUFF1_891 (N3822, N2546);
  buf BUFF1_892 (N3825, N2542);
  buf BUFF1_893 (N3828, N2462);
  buf BUFF1_894 (N3831, N2550);
  buf BUFF1_895 (N3834, N2470);
  buf BUFF1_896 (N3837, N2466);
  buf BUFF1_897 (N3840, N2478);
  buf BUFF1_898 (N3843, N2474);
  buf BUFF1_899 (N3846, N2615);
  buf BUFF1_900 (N3849, N2611);
  buf BUFF1_901 (N3852, N2607);
  buf BUFF1_902 (N3855, N2680);
  buf BUFF1_903 (N3858, N2729);
  buf BUFF1_904 (N3861, N2737);
  buf BUFF1_905 (N3864, N2733);
  buf BUFF1_906 (N3867, N2745);
  buf BUFF1_907 (N3870, N2741);
  buf BUFF1_908 (N3873, N2753);
  buf BUFF1_909 (N3876, N2749);
  buf BUFF1_910 (N3879, N2761);
  buf BUFF1_911 (N3882, N2757);
  or OR2_912 (N3885, N3033, N2419);
  or OR2_913 (N3888, N3032, N2418);
  or OR2_914 (N3891, N3020, N2396);
  nand NAND2_915 (N3953, N3067, N2117);
  not NOT1_916 (N3954, N3067);
  nand NAND2_917 (N3955, N3070, N2537);
  not NOT1_918 (N3956, N3070);
  not NOT1_919 (N3958, N3073);
  not NOT1_920 (N3964, N3080);
  or OR2_921 (N4193, N1649, N3379);
  or OR3_922 (N4303, N1167, N2867, N3130);
  not NOT1_923 (N4308, N3061);
  not NOT1_924 (N4313, N3064);
  nand NAND2_925 (N4326, N2769, N3551);
  nand NAND2_926 (N4327, N2766, N3552);
  nand NAND2_927 (N4333, N2775, N3569);
  nand NAND2_928 (N4334, N2772, N3570);
  nand NAND2_929 (N4411, N2787, N3781);
  nand NAND2_930 (N4412, N2784, N3782);
  nand NAND2_931 (N4463, N3487, N1828);
  not NOT1_932 (N4464, N3487);
  nand NAND2_933 (N4465, N3490, N1829);
  not NOT1_934 (N4466, N3490);
  nand NAND2_935 (N4467, N3493, N2267);
  not NOT1_936 (N4468, N3493);
  nand NAND2_937 (N4469, N3496, N1830);
  not NOT1_938 (N4470, N3496);
  nand NAND2_939 (N4471, N3499, N1833);
  not NOT1_940 (N4472, N3499);
  not NOT1_941 (N4473, N3122);
  not NOT1_942 (N4474, N3126);
  nand NAND2_943 (N4475, N3518, N1840);
  not NOT1_944 (N4476, N3518);
  nand NAND2_945 (N4477, N3521, N1841);
  not NOT1_946 (N4478, N3521);
  nand NAND2_947 (N4479, N3524, N2275);
  not NOT1_948 (N4480, N3524);
  nand NAND2_949 (N4481, N3527, N1842);
  not NOT1_950 (N4482, N3527);
  nand NAND2_951 (N4483, N3530, N1843);
  not NOT1_952 (N4484, N3530);
  not NOT1_953 (N4485, N3155);
  not NOT1_954 (N4486, N3159);
  nand NAND2_955 (N4487, N1721, N3954);
  nand NAND2_956 (N4488, N2235, N3956);
  not NOT1_957 (N4489, N3535);
  nand NAND2_958 (N4490, N3535, N3958);
  not NOT1_959 (N4491, N3539);
  not NOT1_960 (N4492, N3542);
  not NOT1_961 (N4493, N3545);
  not NOT1_962 (N4494, N3548);
  not NOT1_963 (N4495, N3553);
  nand NAND2_964 (N4496, N3553, N3964);
  not NOT1_965 (N4497, N3557);
  not NOT1_966 (N4498, N3560);
  not NOT1_967 (N4499, N3563);
  not NOT1_968 (N4500, N3566);
  not NOT1_969 (N4501, N3571);
  nand NAND2_970 (N4502, N3571, N3167);
  not NOT1_971 (N4503, N3574);
  not NOT1_972 (N4504, N3577);
  not NOT1_973 (N4505, N3580);
  not NOT1_974 (N4506, N3583);
  nand NAND2_975 (N4507, N3598, N1867);
  not NOT1_976 (N4508, N3598);
  nand NAND2_977 (N4509, N3601, N1868);
  not NOT1_978 (N4510, N3601);
  nand NAND2_979 (N4511, N3604, N1869);
  not NOT1_980 (N4512, N3604);
  nand NAND2_981 (N4513, N3607, N1870);
  not NOT1_982 (N4514, N3607);
  nand NAND2_983 (N4515, N3610, N1871);
  not NOT1_984 (N4516, N3610);
  nand NAND2_985 (N4517, N3613, N1872);
  not NOT1_986 (N4518, N3613);
  nand NAND2_987 (N4519, N3616, N1873);
  not NOT1_988 (N4520, N3616);
  nand NAND2_989 (N4521, N3619, N1874);
  not NOT1_990 (N4522, N3619);
  nand NAND2_991 (N4523, N3622, N1875);
  not NOT1_992 (N4524, N3622);
  nand NAND2_993 (N4525, N3631, N1876);
  not NOT1_994 (N4526, N3631);
  nand NAND2_995 (N4527, N3634, N1877);
  not NOT1_996 (N4528, N3634);
  nand NAND2_997 (N4529, N3637, N1878);
  not NOT1_998 (N4530, N3637);
  nand NAND2_999 (N4531, N3640, N1879);
  not NOT1_1000 (N4532, N3640);
  nand NAND2_1001 (N4533, N3643, N1880);
  not NOT1_1002 (N4534, N3643);
  nand NAND2_1003 (N4535, N3646, N1881);
  not NOT1_1004 (N4536, N3646);
  nand NAND2_1005 (N4537, N3649, N1882);
  not NOT1_1006 (N4538, N3649);
  nand NAND2_1007 (N4539, N3652, N1883);
  not NOT1_1008 (N4540, N3652);
  nand NAND2_1009 (N4541, N3655, N1884);
  not NOT1_1010 (N4542, N3655);
  not NOT1_1011 (N4543, N3658);
  and AND2_1012 (N4544, N806, N3293);
  and AND2_1013 (N4545, N800, N3287);
  and AND2_1014 (N4549, N794, N3281);
  and AND2_1015 (N4555, N3273, N786);
  and AND2_1016 (N4562, N780, N3267);
  and AND2_1017 (N4563, N774, N3355);
  and AND2_1018 (N4566, N768, N3349);
  and AND2_1019 (N4570, N762, N3343);
  not NOT1_1020 (N4575, N3661);
  and AND2_1021 (N4576, N806, N3293);
  and AND2_1022 (N4577, N800, N3287);
  and AND2_1023 (N4581, N794, N3281);
  and AND2_1024 (N4586, N786, N3273);
  and AND2_1025 (N4592, N780, N3267);
  and AND2_1026 (N4593, N774, N3355);
  and AND2_1027 (N4597, N768, N3349);
  and AND2_1028 (N4603, N762, N3343);
  not NOT1_1029 (N4610, N3664);
  not NOT1_1030 (N4611, N3667);
  not NOT1_1031 (N4612, N3670);
  not NOT1_1032 (N4613, N3673);
  not NOT1_1033 (N4614, N3676);
  not NOT1_1034 (N4615, N3679);
  not NOT1_1035 (N4616, N3682);
  not NOT1_1036 (N4617, N3685);
  not NOT1_1037 (N4618, N3688);
  not NOT1_1038 (N4619, N3691);
  not NOT1_1039 (N4620, N3694);
  not NOT1_1040 (N4621, N3697);
  not NOT1_1041 (N4622, N3700);
  not NOT1_1042 (N4623, N3703);
  not NOT1_1043 (N4624, N3706);
  not NOT1_1044 (N4625, N3709);
  not NOT1_1045 (N4626, N3712);
  not NOT1_1046 (N4627, N3715);
  not NOT1_1047 (N4628, N3718);
  not NOT1_1048 (N4629, N3721);
  and AND2_1049 (N4630, N3448, N2704);
  not NOT1_1050 (N4631, N3724);
  and AND2_1051 (N4632, N3444, N2700);
  not NOT1_1052 (N4633, N3727);
  and AND2_1053 (N4634, N3440, N2696);
  and AND2_1054 (N4635, N3436, N2692);
  not NOT1_1055 (N4636, N3730);
  and AND2_1056 (N4637, N3432, N2688);
  and AND2_1057 (N4638, N3428, N3311);
  and AND2_1058 (N4639, N3424, N3307);
  and AND2_1059 (N4640, N3420, N3303);
  and AND2_1060 (N4641, N3416, N3299);
  not NOT1_1061 (N4642, N3733);
  not NOT1_1062 (N4643, N3736);
  not NOT1_1063 (N4644, N3739);
  not NOT1_1064 (N4645, N3742);
  not NOT1_1065 (N4646, N3745);
  not NOT1_1066 (N4647, N3748);
  not NOT1_1067 (N4648, N3751);
  not NOT1_1068 (N4649, N3754);
  not NOT1_1069 (N4650, N3757);
  not NOT1_1070 (N4651, N3760);
  not NOT1_1071 (N4652, N3763);
  not NOT1_1072 (N4653, N3375);
  and AND2_1073 (N4656, N865, N3410);
  and AND2_1074 (N4657, N859, N3404);
  and AND2_1075 (N4661, N853, N3398);
  and AND2_1076 (N4667, N3390, N845);
  and AND2_1077 (N4674, N839, N3384);
  and AND2_1078 (N4675, N833, N3334);
  and AND2_1079 (N4678, N827, N3328);
  and AND2_1080 (N4682, N821, N3322);
  and AND2_1081 (N4687, N814, N3315);
  not NOT1_1082 (N4693, N3766);
  nand NAND2_1083 (N4694, N3766, N3380);
  not NOT1_1084 (N4695, N3769);
  not NOT1_1085 (N4696, N3772);
  not NOT1_1086 (N4697, N3775);
  not NOT1_1087 (N4698, N3778);
  not NOT1_1088 (N4699, N3783);
  not NOT1_1089 (N4700, N3786);
  and AND2_1090 (N4701, N865, N3410);
  and AND2_1091 (N4702, N859, N3404);
  and AND2_1092 (N4706, N853, N3398);
  and AND2_1093 (N4711, N845, N3390);
  and AND2_1094 (N4717, N839, N3384);
  and AND2_1095 (N4718, N833, N3334);
  and AND2_1096 (N4722, N827, N3328);
  and AND2_1097 (N4728, N821, N3322);
  and AND2_1098 (N4735, N814, N3315);
  not NOT1_1099 (N4743, N3789);
  not NOT1_1100 (N4744, N3792);
  not NOT1_1101 (N4745, N3807);
  nand NAND2_1102 (N4746, N3807, N3452);
  not NOT1_1103 (N4747, N3810);
  not NOT1_1104 (N4748, N3813);
  not NOT1_1105 (N4749, N3816);
  not NOT1_1106 (N4750, N3819);
  nand NAND2_1107 (N4751, N3819, N3453);
  not NOT1_1108 (N4752, N3822);
  not NOT1_1109 (N4753, N3825);
  not NOT1_1110 (N4754, N3828);
  not NOT1_1111 (N4755, N3831);
  and AND2_1112 (N4756, N3482, N3263);
  and AND2_1113 (N4757, N3478, N3259);
  and AND2_1114 (N4758, N3474, N3255);
  and AND2_1115 (N4759, N3470, N3251);
  and AND2_1116 (N4760, N3466, N3247);
  not NOT1_1117 (N4761, N3846);
  and AND2_1118 (N4762, N3462, N2615);
  not NOT1_1119 (N4763, N3849);
  and AND2_1120 (N4764, N3458, N2611);
  not NOT1_1121 (N4765, N3852);
  and AND2_1122 (N4766, N3454, N2607);
  and AND2_1123 (N4767, N2680, N3381);
  not NOT1_1124 (N4768, N3855);
  and AND2_1125 (N4769, N3340, N695);
  not NOT1_1126 (N4775, N3858);
  nand NAND2_1127 (N4776, N3858, N3486);
  not NOT1_1128 (N4777, N3861);
  not NOT1_1129 (N4778, N3864);
  not NOT1_1130 (N4779, N3867);
  not NOT1_1131 (N4780, N3870);
  not NOT1_1132 (N4781, N3885);
  not NOT1_1133 (N4782, N3888);
  not NOT1_1134 (N4783, N3891);
  or OR2_1135 (N4784, N3131, N3134);
  not NOT1_1136 (N4789, N3502);
  not NOT1_1137 (N4790, N3131);
  not NOT1_1138 (N4793, N3507);
  not NOT1_1139 (N4794, N3510);
  not NOT1_1140 (N4795, N3515);
  buf BUFF1_1141 (N4796, N3114);
  not NOT1_1142 (N4799, N3586);
  not NOT1_1143 (N4800, N3589);
  not NOT1_1144 (N4801, N3592);
  not NOT1_1145 (N4802, N3595);
  nand NAND2_1146 (N4803, N4326, N4327);
  nand NAND2_1147 (N4806, N4333, N4334);
  not NOT1_1148 (N4809, N3625);
  buf BUFF1_1149 (N4810, N3178);
  not NOT1_1150 (N4813, N3628);
  buf BUFF1_1151 (N4814, N3202);
  buf BUFF1_1152 (N4817, N3221);
  buf BUFF1_1153 (N4820, N3293);
  buf BUFF1_1154 (N4823, N3287);
  buf BUFF1_1155 (N4826, N3281);
  buf BUFF1_1156 (N4829, N3273);
  buf BUFF1_1157 (N4832, N3267);
  buf BUFF1_1158 (N4835, N3355);
  buf BUFF1_1159 (N4838, N3349);
  buf BUFF1_1160 (N4841, N3343);
  nor NOR2_1161 (N4844, N3273, N786);
  buf BUFF1_1162 (N4847, N3293);
  buf BUFF1_1163 (N4850, N3287);
  buf BUFF1_1164 (N4853, N3281);
  buf BUFF1_1165 (N4856, N3267);
  buf BUFF1_1166 (N4859, N3355);
  buf BUFF1_1167 (N4862, N3349);
  buf BUFF1_1168 (N4865, N3343);
  buf BUFF1_1169 (N4868, N3273);
  nor NOR2_1170 (N4871, N786, N3273);
  buf BUFF1_1171 (N4874, N3448);
  buf BUFF1_1172 (N4877, N3444);
  buf BUFF1_1173 (N4880, N3440);
  buf BUFF1_1174 (N4883, N3432);
  buf BUFF1_1175 (N4886, N3428);
  buf BUFF1_1176 (N4889, N3311);
  buf BUFF1_1177 (N4892, N3424);
  buf BUFF1_1178 (N4895, N3307);
  buf BUFF1_1179 (N4898, N3420);
  buf BUFF1_1180 (N4901, N3303);
  buf BUFF1_1181 (N4904, N3436);
  buf BUFF1_1182 (N4907, N3416);
  buf BUFF1_1183 (N4910, N3299);
  buf BUFF1_1184 (N4913, N3410);
  buf BUFF1_1185 (N4916, N3404);
  buf BUFF1_1186 (N4919, N3398);
  buf BUFF1_1187 (N4922, N3390);
  buf BUFF1_1188 (N4925, N3384);
  buf BUFF1_1189 (N4928, N3334);
  buf BUFF1_1190 (N4931, N3328);
  buf BUFF1_1191 (N4934, N3322);
  buf BUFF1_1192 (N4937, N3315);
  nor NOR2_1193 (N4940, N3390, N845);
  buf BUFF1_1194 (N4943, N3315);
  buf BUFF1_1195 (N4946, N3328);
  buf BUFF1_1196 (N4949, N3322);
  buf BUFF1_1197 (N4952, N3384);
  buf BUFF1_1198 (N4955, N3334);
  buf BUFF1_1199 (N4958, N3398);
  buf BUFF1_1200 (N4961, N3390);
  buf BUFF1_1201 (N4964, N3410);
  buf BUFF1_1202 (N4967, N3404);
  buf BUFF1_1203 (N4970, N3340);
  buf BUFF1_1204 (N4973, N3349);
  buf BUFF1_1205 (N4976, N3343);
  buf BUFF1_1206 (N4979, N3267);
  buf BUFF1_1207 (N4982, N3355);
  buf BUFF1_1208 (N4985, N3281);
  buf BUFF1_1209 (N4988, N3273);
  buf BUFF1_1210 (N4991, N3293);
  buf BUFF1_1211 (N4994, N3287);
  nand NAND2_1212 (N4997, N4411, N4412);
  buf BUFF1_1213 (N5000, N3410);
  buf BUFF1_1214 (N5003, N3404);
  buf BUFF1_1215 (N5006, N3398);
  buf BUFF1_1216 (N5009, N3384);
  buf BUFF1_1217 (N5012, N3334);
  buf BUFF1_1218 (N5015, N3328);
  buf BUFF1_1219 (N5018, N3322);
  buf BUFF1_1220 (N5021, N3390);
  buf BUFF1_1221 (N5024, N3315);
  nor NOR2_1222 (N5027, N845, N3390);
  nor NOR2_1223 (N5030, N814, N3315);
  buf BUFF1_1224 (N5033, N3299);
  buf BUFF1_1225 (N5036, N3307);
  buf BUFF1_1226 (N5039, N3303);
  buf BUFF1_1227 (N5042, N3311);
  not NOT1_1228 (N5045, N3795);
  not NOT1_1229 (N5046, N3798);
  not NOT1_1230 (N5047, N3801);
  not NOT1_1231 (N5048, N3804);
  buf BUFF1_1232 (N5049, N3247);
  buf BUFF1_1233 (N5052, N3255);
  buf BUFF1_1234 (N5055, N3251);
  buf BUFF1_1235 (N5058, N3263);
  buf BUFF1_1236 (N5061, N3259);
  not NOT1_1237 (N5064, N3834);
  not NOT1_1238 (N5065, N3837);
  not NOT1_1239 (N5066, N3840);
  not NOT1_1240 (N5067, N3843);
  buf BUFF1_1241 (N5068, N3482);
  buf BUFF1_1242 (N5071, N3263);
  buf BUFF1_1243 (N5074, N3478);
  buf BUFF1_1244 (N5077, N3259);
  buf BUFF1_1245 (N5080, N3474);
  buf BUFF1_1246 (N5083, N3255);
  buf BUFF1_1247 (N5086, N3466);
  buf BUFF1_1248 (N5089, N3247);
  buf BUFF1_1249 (N5092, N3462);
  buf BUFF1_1250 (N5095, N3458);
  buf BUFF1_1251 (N5098, N3454);
  buf BUFF1_1252 (N5101, N3470);
  buf BUFF1_1253 (N5104, N3251);
  buf BUFF1_1254 (N5107, N3381);
  not NOT1_1255 (N5110, N3873);
  not NOT1_1256 (N5111, N3876);
  not NOT1_1257 (N5112, N3879);
  not NOT1_1258 (N5113, N3882);
  buf BUFF1_1259 (N5114, N3458);
  buf BUFF1_1260 (N5117, N3454);
  buf BUFF1_1261 (N5120, N3466);
  buf BUFF1_1262 (N5123, N3462);
  buf BUFF1_1263 (N5126, N3474);
  buf BUFF1_1264 (N5129, N3470);
  buf BUFF1_1265 (N5132, N3482);
  buf BUFF1_1266 (N5135, N3478);
  buf BUFF1_1267 (N5138, N3416);
  buf BUFF1_1268 (N5141, N3424);
  buf BUFF1_1269 (N5144, N3420);
  buf BUFF1_1270 (N5147, N3432);
  buf BUFF1_1271 (N5150, N3428);
  buf BUFF1_1272 (N5153, N3440);
  buf BUFF1_1273 (N5156, N3436);
  buf BUFF1_1274 (N5159, N3448);
  buf BUFF1_1275 (N5162, N3444);
  nand NAND2_1276 (N5165, N4486, N4485);
  nand NAND2_1277 (N5166, N4474, N4473);
  nand NAND2_1278 (N5167, N1290, N4464);
  nand NAND2_1279 (N5168, N1293, N4466);
  nand NAND2_1280 (N5169, N2074, N4468);
  nand NAND2_1281 (N5170, N1296, N4470);
  nand NAND2_1282 (N5171, N1302, N4472);
  nand NAND2_1283 (N5172, N1314, N4476);
  nand NAND2_1284 (N5173, N1317, N4478);
  nand NAND2_1285 (N5174, N2081, N4480);
  nand NAND2_1286 (N5175, N1320, N4482);
  nand NAND2_1287 (N5176, N1323, N4484);
  nand NAND2_1288 (N5177, N3953, N4487);
  nand NAND2_1289 (N5178, N3955, N4488);
  nand NAND2_1290 (N5179, N3073, N4489);
  nand NAND2_1291 (N5180, N3542, N4491);
  nand NAND2_1292 (N5181, N3539, N4492);
  nand NAND2_1293 (N5182, N3548, N4493);
  nand NAND2_1294 (N5183, N3545, N4494);
  nand NAND2_1295 (N5184, N3080, N4495);
  nand NAND2_1296 (N5185, N3560, N4497);
  nand NAND2_1297 (N5186, N3557, N4498);
  nand NAND2_1298 (N5187, N3566, N4499);
  nand NAND2_1299 (N5188, N3563, N4500);
  nand NAND2_1300 (N5189, N2778, N4501);
  nand NAND2_1301 (N5190, N3577, N4503);
  nand NAND2_1302 (N5191, N3574, N4504);
  nand NAND2_1303 (N5192, N3583, N4505);
  nand NAND2_1304 (N5193, N3580, N4506);
  nand NAND2_1305 (N5196, N1326, N4508);
  nand NAND2_1306 (N5197, N1329, N4510);
  nand NAND2_1307 (N5198, N1332, N4512);
  nand NAND2_1308 (N5199, N1335, N4514);
  nand NAND2_1309 (N5200, N1338, N4516);
  nand NAND2_1310 (N5201, N1341, N4518);
  nand NAND2_1311 (N5202, N1344, N4520);
  nand NAND2_1312 (N5203, N1347, N4522);
  nand NAND2_1313 (N5204, N1350, N4524);
  nand NAND2_1314 (N5205, N1353, N4526);
  nand NAND2_1315 (N5206, N1356, N4528);
  nand NAND2_1316 (N5207, N1359, N4530);
  nand NAND2_1317 (N5208, N1362, N4532);
  nand NAND2_1318 (N5209, N1365, N4534);
  nand NAND2_1319 (N5210, N1368, N4536);
  nand NAND2_1320 (N5211, N1371, N4538);
  nand NAND2_1321 (N5212, N1374, N4540);
  nand NAND2_1322 (N5213, N1377, N4542);
  nand NAND2_1323 (N5283, N3670, N4611);
  nand NAND2_1324 (N5284, N3667, N4612);
  nand NAND2_1325 (N5285, N3676, N4613);
  nand NAND2_1326 (N5286, N3673, N4614);
  nand NAND2_1327 (N5287, N3682, N4615);
  nand NAND2_1328 (N5288, N3679, N4616);
  nand NAND2_1329 (N5289, N3688, N4617);
  nand NAND2_1330 (N5290, N3685, N4618);
  nand NAND2_1331 (N5291, N3694, N4619);
  nand NAND2_1332 (N5292, N3691, N4620);
  nand NAND2_1333 (N5293, N3700, N4621);
  nand NAND2_1334 (N5294, N3697, N4622);
  nand NAND2_1335 (N5295, N3706, N4623);
  nand NAND2_1336 (N5296, N3703, N4624);
  nand NAND2_1337 (N5297, N3712, N4625);
  nand NAND2_1338 (N5298, N3709, N4626);
  nand NAND2_1339 (N5299, N3718, N4627);
  nand NAND2_1340 (N5300, N3715, N4628);
  nand NAND2_1341 (N5314, N3739, N4643);
  nand NAND2_1342 (N5315, N3736, N4644);
  nand NAND2_1343 (N5316, N3745, N4645);
  nand NAND2_1344 (N5317, N3742, N4646);
  nand NAND2_1345 (N5318, N3751, N4647);
  nand NAND2_1346 (N5319, N3748, N4648);
  nand NAND2_1347 (N5320, N3757, N4649);
  nand NAND2_1348 (N5321, N3754, N4650);
  nand NAND2_1349 (N5322, N3763, N4651);
  nand NAND2_1350 (N5323, N3760, N4652);
  not NOT1_1351 (N5324, N4193);
  nand NAND2_1352 (N5363, N2781, N4693);
  nand NAND2_1353 (N5364, N3772, N4695);
  nand NAND2_1354 (N5365, N3769, N4696);
  nand NAND2_1355 (N5366, N3778, N4697);
  nand NAND2_1356 (N5367, N3775, N4698);
  nand NAND2_1357 (N5425, N2790, N4745);
  nand NAND2_1358 (N5426, N3813, N4747);
  nand NAND2_1359 (N5427, N3810, N4748);
  nand NAND2_1360 (N5429, N2793, N4750);
  nand NAND2_1361 (N5430, N3825, N4752);
  nand NAND2_1362 (N5431, N3822, N4753);
  nand NAND2_1363 (N5432, N3831, N4754);
  nand NAND2_1364 (N5433, N3828, N4755);
  nand NAND2_1365 (N5451, N2796, N4775);
  nand NAND2_1366 (N5452, N3864, N4777);
  nand NAND2_1367 (N5453, N3861, N4778);
  nand NAND2_1368 (N5454, N3870, N4779);
  nand NAND2_1369 (N5455, N3867, N4780);
  nand NAND2_1370 (N5456, N3888, N4781);
  nand NAND2_1371 (N5457, N3885, N4782);
  not NOT1_1372 (N5469, N4303);
  nand NAND2_1373 (N5474, N3589, N4799);
  nand NAND2_1374 (N5475, N3586, N4800);
  nand NAND2_1375 (N5476, N3595, N4801);
  nand NAND2_1376 (N5477, N3592, N4802);
  nand NAND2_1377 (N5571, N3798, N5045);
  nand NAND2_1378 (N5572, N3795, N5046);
  nand NAND2_1379 (N5573, N3804, N5047);
  nand NAND2_1380 (N5574, N3801, N5048);
  nand NAND2_1381 (N5584, N3837, N5064);
  nand NAND2_1382 (N5585, N3834, N5065);
  nand NAND2_1383 (N5586, N3843, N5066);
  nand NAND2_1384 (N5587, N3840, N5067);
  nand NAND2_1385 (N5602, N3876, N5110);
  nand NAND2_1386 (N5603, N3873, N5111);
  nand NAND2_1387 (N5604, N3882, N5112);
  nand NAND2_1388 (N5605, N3879, N5113);
  nand NAND2_1389 (N5631, N5324, N4653);
  nand NAND2_1390 (N5632, N4463, N5167);
  nand NAND2_1391 (N5640, N4465, N5168);
  nand NAND2_1392 (N5654, N4467, N5169);
  nand NAND2_1393 (N5670, N4469, N5170);
  nand NAND2_1394 (N5683, N4471, N5171);
  nand NAND2_1395 (N5690, N4475, N5172);
  nand NAND2_1396 (N5697, N4477, N5173);
  nand NAND2_1397 (N5707, N4479, N5174);
  nand NAND2_1398 (N5718, N4481, N5175);
  nand NAND2_1399 (N5728, N4483, N5176);
  not NOT1_1400 (N5735, N5177);
  nand NAND2_1401 (N5736, N5179, N4490);
  nand NAND2_1402 (N5740, N5180, N5181);
  nand NAND2_1403 (N5744, N5182, N5183);
  nand NAND2_1404 (N5747, N5184, N4496);
  nand NAND2_1405 (N5751, N5185, N5186);
  nand NAND2_1406 (N5755, N5187, N5188);
  nand NAND2_1407 (N5758, N5189, N4502);
  nand NAND2_1408 (N5762, N5190, N5191);
  nand NAND2_1409 (N5766, N5192, N5193);
  not NOT1_1410 (N5769, N4803);
  not NOT1_1411 (N5770, N4806);
  nand NAND2_1412 (N5771, N4507, N5196);
  nand NAND2_1413 (N5778, N4509, N5197);
  nand NAND2_1414 (N5789, N4511, N5198);
  nand NAND2_1415 (N5799, N4513, N5199);
  nand NAND2_1416 (N5807, N4515, N5200);
  nand NAND2_1417 (N5821, N4517, N5201);
  nand NAND2_1418 (N5837, N4519, N5202);
  nand NAND2_1419 (N5850, N4521, N5203);
  nand NAND2_1420 (N5856, N4523, N5204);
  nand NAND2_1421 (N5863, N4525, N5205);
  nand NAND2_1422 (N5870, N4527, N5206);
  nand NAND2_1423 (N5881, N4529, N5207);
  nand NAND2_1424 (N5892, N4531, N5208);
  nand NAND2_1425 (N5898, N4533, N5209);
  nand NAND2_1426 (N5905, N4535, N5210);
  nand NAND2_1427 (N5915, N4537, N5211);
  nand NAND2_1428 (N5926, N4539, N5212);
  nand NAND2_1429 (N5936, N4541, N5213);
  not NOT1_1430 (N5943, N4817);
  nand NAND2_1431 (N5944, N4820, N1931);
  not NOT1_1432 (N5945, N4820);
  nand NAND2_1433 (N5946, N4823, N1932);
  not NOT1_1434 (N5947, N4823);
  nand NAND2_1435 (N5948, N4826, N1933);
  not NOT1_1436 (N5949, N4826);
  nand NAND2_1437 (N5950, N4829, N1934);
  not NOT1_1438 (N5951, N4829);
  nand NAND2_1439 (N5952, N4832, N1935);
  not NOT1_1440 (N5953, N4832);
  nand NAND2_1441 (N5954, N4835, N1936);
  not NOT1_1442 (N5955, N4835);
  nand NAND2_1443 (N5956, N4838, N1937);
  not NOT1_1444 (N5957, N4838);
  nand NAND2_1445 (N5958, N4841, N1938);
  not NOT1_1446 (N5959, N4841);
  and AND2_1447 (N5960, N2674, N4769);
  not NOT1_1448 (N5966, N4844);
  nand NAND2_1449 (N5967, N4847, N1939);
  not NOT1_1450 (N5968, N4847);
  nand NAND2_1451 (N5969, N4850, N1940);
  not NOT1_1452 (N5970, N4850);
  nand NAND2_1453 (N5971, N4853, N1941);
  not NOT1_1454 (N5972, N4853);
  nand NAND2_1455 (N5973, N4856, N1942);
  not NOT1_1456 (N5974, N4856);
  nand NAND2_1457 (N5975, N4859, N1943);
  not NOT1_1458 (N5976, N4859);
  nand NAND2_1459 (N5977, N4862, N1944);
  not NOT1_1460 (N5978, N4862);
  nand NAND2_1461 (N5979, N4865, N1945);
  not NOT1_1462 (N5980, N4865);
  and AND2_1463 (N5981, N2674, N4769);
  nand NAND2_1464 (N5989, N4868, N1946);
  not NOT1_1465 (N5990, N4868);
  nand NAND2_1466 (N5991, N5283, N5284);
  nand NAND2_1467 (N5996, N5285, N5286);
  nand NAND2_1468 (N6000, N5287, N5288);
  nand NAND2_1469 (N6003, N5289, N5290);
  nand NAND2_1470 (N6009, N5291, N5292);
  nand NAND2_1471 (N6014, N5293, N5294);
  nand NAND2_1472 (N6018, N5295, N5296);
  nand NAND2_1473 (N6021, N5297, N5298);
  nand NAND2_1474 (N6022, N5299, N5300);
  not NOT1_1475 (N6023, N4874);
  nand NAND2_1476 (N6024, N4874, N4629);
  not NOT1_1477 (N6025, N4877);
  nand NAND2_1478 (N6026, N4877, N4631);
  not NOT1_1479 (N6027, N4880);
  nand NAND2_1480 (N6028, N4880, N4633);
  not NOT1_1481 (N6029, N4883);
  nand NAND2_1482 (N6030, N4883, N4636);
  not NOT1_1483 (N6031, N4886);
  not NOT1_1484 (N6032, N4889);
  not NOT1_1485 (N6033, N4892);
  not NOT1_1486 (N6034, N4895);
  not NOT1_1487 (N6035, N4898);
  not NOT1_1488 (N6036, N4901);
  not NOT1_1489 (N6037, N4904);
  nand NAND2_1490 (N6038, N4904, N4642);
  not NOT1_1491 (N6039, N4907);
  not NOT1_1492 (N6040, N4910);
  nand NAND2_1493 (N6041, N5314, N5315);
  nand NAND2_1494 (N6047, N5316, N5317);
  nand NAND2_1495 (N6052, N5318, N5319);
  nand NAND2_1496 (N6056, N5320, N5321);
  nand NAND2_1497 (N6059, N5322, N5323);
  nand NAND2_1498 (N6060, N4913, N1968);
  not NOT1_1499 (N6061, N4913);
  nand NAND2_1500 (N6062, N4916, N1969);
  not NOT1_1501 (N6063, N4916);
  nand NAND2_1502 (N6064, N4919, N1970);
  not NOT1_1503 (N6065, N4919);
  nand NAND2_1504 (N6066, N4922, N1971);
  not NOT1_1505 (N6067, N4922);
  nand NAND2_1506 (N6068, N4925, N1972);
  not NOT1_1507 (N6069, N4925);
  nand NAND2_1508 (N6070, N4928, N1973);
  not NOT1_1509 (N6071, N4928);
  nand NAND2_1510 (N6072, N4931, N1974);
  not NOT1_1511 (N6073, N4931);
  nand NAND2_1512 (N6074, N4934, N1975);
  not NOT1_1513 (N6075, N4934);
  nand NAND2_1514 (N6076, N4937, N1976);
  not NOT1_1515 (N6077, N4937);
  not NOT1_1516 (N6078, N4940);
  nand NAND2_1517 (N6079, N5363, N4694);
  nand NAND2_1518 (N6083, N5364, N5365);
  nand NAND2_1519 (N6087, N5366, N5367);
  not NOT1_1520 (N6090, N4943);
  nand NAND2_1521 (N6091, N4943, N4699);
  not NOT1_1522 (N6092, N4946);
  not NOT1_1523 (N6093, N4949);
  not NOT1_1524 (N6094, N4952);
  not NOT1_1525 (N6095, N4955);
  not NOT1_1526 (N6096, N4970);
  nand NAND2_1527 (N6097, N4970, N4700);
  not NOT1_1528 (N6098, N4973);
  not NOT1_1529 (N6099, N4976);
  not NOT1_1530 (N6100, N4979);
  not NOT1_1531 (N6101, N4982);
  not NOT1_1532 (N6102, N4997);
  nand NAND2_1533 (N6103, N5000, N2015);
  not NOT1_1534 (N6104, N5000);
  nand NAND2_1535 (N6105, N5003, N2016);
  not NOT1_1536 (N6106, N5003);
  nand NAND2_1537 (N6107, N5006, N2017);
  not NOT1_1538 (N6108, N5006);
  nand NAND2_1539 (N6109, N5009, N2018);
  not NOT1_1540 (N6110, N5009);
  nand NAND2_1541 (N6111, N5012, N2019);
  not NOT1_1542 (N6112, N5012);
  nand NAND2_1543 (N6113, N5015, N2020);
  not NOT1_1544 (N6114, N5015);
  nand NAND2_1545 (N6115, N5018, N2021);
  not NOT1_1546 (N6116, N5018);
  nand NAND2_1547 (N6117, N5021, N2022);
  not NOT1_1548 (N6118, N5021);
  nand NAND2_1549 (N6119, N5024, N2023);
  not NOT1_1550 (N6120, N5024);
  not NOT1_1551 (N6121, N5033);
  nand NAND2_1552 (N6122, N5033, N4743);
  not NOT1_1553 (N6123, N5036);
  not NOT1_1554 (N6124, N5039);
  nand NAND2_1555 (N6125, N5042, N4744);
  not NOT1_1556 (N6126, N5042);
  nand NAND2_1557 (N6127, N5425, N4746);
  nand NAND2_1558 (N6131, N5426, N5427);
  not NOT1_1559 (N6135, N5049);
  nand NAND2_1560 (N6136, N5049, N4749);
  nand NAND2_1561 (N6137, N5429, N4751);
  nand NAND2_1562 (N6141, N5430, N5431);
  nand NAND2_1563 (N6145, N5432, N5433);
  not NOT1_1564 (N6148, N5068);
  not NOT1_1565 (N6149, N5071);
  not NOT1_1566 (N6150, N5074);
  not NOT1_1567 (N6151, N5077);
  not NOT1_1568 (N6152, N5080);
  not NOT1_1569 (N6153, N5083);
  not NOT1_1570 (N6154, N5086);
  not NOT1_1571 (N6155, N5089);
  not NOT1_1572 (N6156, N5092);
  nand NAND2_1573 (N6157, N5092, N4761);
  not NOT1_1574 (N6158, N5095);
  nand NAND2_1575 (N6159, N5095, N4763);
  not NOT1_1576 (N6160, N5098);
  nand NAND2_1577 (N6161, N5098, N4765);
  not NOT1_1578 (N6162, N5101);
  not NOT1_1579 (N6163, N5104);
  nand NAND2_1580 (N6164, N5107, N4768);
  not NOT1_1581 (N6165, N5107);
  nand NAND2_1582 (N6166, N5451, N4776);
  nand NAND2_1583 (N6170, N5452, N5453);
  nand NAND2_1584 (N6174, N5454, N5455);
  nand NAND2_1585 (N6177, N5456, N5457);
  not NOT1_1586 (N6181, N5114);
  not NOT1_1587 (N6182, N5117);
  not NOT1_1588 (N6183, N5120);
  not NOT1_1589 (N6184, N5123);
  not NOT1_1590 (N6185, N5138);
  nand NAND2_1591 (N6186, N5138, N4783);
  not NOT1_1592 (N6187, N5141);
  not NOT1_1593 (N6188, N5144);
  not NOT1_1594 (N6189, N5147);
  not NOT1_1595 (N6190, N5150);
  not NOT1_1596 (N6191, N4784);
  nand NAND2_1597 (N6192, N4784, N2230);
  not NOT1_1598 (N6193, N4790);
  nand NAND2_1599 (N6194, N4790, N2765);
  not NOT1_1600 (N6195, N4796);
  nand NAND2_1601 (N6196, N5476, N5477);
  nand NAND2_1602 (N6199, N5474, N5475);
  not NOT1_1603 (N6202, N4810);
  not NOT1_1604 (N6203, N4814);
  buf BUFF1_1605 (N6204, N4769);
  buf BUFF1_1606 (N6207, N4555);
  buf BUFF1_1607 (N6210, N4769);
  not NOT1_1608 (N6213, N4871);
  buf BUFF1_1609 (N6214, N4586);
  nor NOR2_1610 (N6217, N2674, N4769);
  buf BUFF1_1611 (N6220, N4667);
  not NOT1_1612 (N6223, N4958);
  not NOT1_1613 (N6224, N4961);
  not NOT1_1614 (N6225, N4964);
  not NOT1_1615 (N6226, N4967);
  not NOT1_1616 (N6227, N4985);
  not NOT1_1617 (N6228, N4988);
  not NOT1_1618 (N6229, N4991);
  not NOT1_1619 (N6230, N4994);
  not NOT1_1620 (N6231, N5027);
  buf BUFF1_1621 (N6232, N4711);
  not NOT1_1622 (N6235, N5030);
  buf BUFF1_1623 (N6236, N4735);
  not NOT1_1624 (N6239, N5052);
  not NOT1_1625 (N6240, N5055);
  not NOT1_1626 (N6241, N5058);
  not NOT1_1627 (N6242, N5061);
  nand NAND2_1628 (N6243, N5573, N5574);
  nand NAND2_1629 (N6246, N5571, N5572);
  nand NAND2_1630 (N6249, N5586, N5587);
  nand NAND2_1631 (N6252, N5584, N5585);
  not NOT1_1632 (N6255, N5126);
  not NOT1_1633 (N6256, N5129);
  not NOT1_1634 (N6257, N5132);
  not NOT1_1635 (N6258, N5135);
  not NOT1_1636 (N6259, N5153);
  not NOT1_1637 (N6260, N5156);
  not NOT1_1638 (N6261, N5159);
  not NOT1_1639 (N6262, N5162);
  nand NAND2_1640 (N6263, N5604, N5605);
  nand NAND2_1641 (N6266, N5602, N5603);
  nand NAND2_1642 (N6540, N1380, N5945);
  nand NAND2_1643 (N6541, N1383, N5947);
  nand NAND2_1644 (N6542, N1386, N5949);
  nand NAND2_1645 (N6543, N1389, N5951);
  nand NAND2_1646 (N6544, N1392, N5953);
  nand NAND2_1647 (N6545, N1395, N5955);
  nand NAND2_1648 (N6546, N1398, N5957);
  nand NAND2_1649 (N6547, N1401, N5959);
  nand NAND2_1650 (N6555, N1404, N5968);
  nand NAND2_1651 (N6556, N1407, N5970);
  nand NAND2_1652 (N6557, N1410, N5972);
  nand NAND2_1653 (N6558, N1413, N5974);
  nand NAND2_1654 (N6559, N1416, N5976);
  nand NAND2_1655 (N6560, N1419, N5978);
  nand NAND2_1656 (N6561, N1422, N5980);
  nand NAND2_1657 (N6569, N1425, N5990);
  nand NAND2_1658 (N6594, N3721, N6023);
  nand NAND2_1659 (N6595, N3724, N6025);
  nand NAND2_1660 (N6596, N3727, N6027);
  nand NAND2_1661 (N6597, N3730, N6029);
  nand NAND2_1662 (N6598, N4889, N6031);
  nand NAND2_1663 (N6599, N4886, N6032);
  nand NAND2_1664 (N6600, N4895, N6033);
  nand NAND2_1665 (N6601, N4892, N6034);
  nand NAND2_1666 (N6602, N4901, N6035);
  nand NAND2_1667 (N6603, N4898, N6036);
  nand NAND2_1668 (N6604, N3733, N6037);
  nand NAND2_1669 (N6605, N4910, N6039);
  nand NAND2_1670 (N6606, N4907, N6040);
  nand NAND2_1671 (N6621, N1434, N6061);
  nand NAND2_1672 (N6622, N1437, N6063);
  nand NAND2_1673 (N6623, N1440, N6065);
  nand NAND2_1674 (N6624, N1443, N6067);
  nand NAND2_1675 (N6625, N1446, N6069);
  nand NAND2_1676 (N6626, N1449, N6071);
  nand NAND2_1677 (N6627, N1452, N6073);
  nand NAND2_1678 (N6628, N1455, N6075);
  nand NAND2_1679 (N6629, N1458, N6077);
  nand NAND2_1680 (N6639, N3783, N6090);
  nand NAND2_1681 (N6640, N4949, N6092);
  nand NAND2_1682 (N6641, N4946, N6093);
  nand NAND2_1683 (N6642, N4955, N6094);
  nand NAND2_1684 (N6643, N4952, N6095);
  nand NAND2_1685 (N6644, N3786, N6096);
  nand NAND2_1686 (N6645, N4976, N6098);
  nand NAND2_1687 (N6646, N4973, N6099);
  nand NAND2_1688 (N6647, N4982, N6100);
  nand NAND2_1689 (N6648, N4979, N6101);
  nand NAND2_1690 (N6649, N1461, N6104);
  nand NAND2_1691 (N6650, N1464, N6106);
  nand NAND2_1692 (N6651, N1467, N6108);
  nand NAND2_1693 (N6652, N1470, N6110);
  nand NAND2_1694 (N6653, N1473, N6112);
  nand NAND2_1695 (N6654, N1476, N6114);
  nand NAND2_1696 (N6655, N1479, N6116);
  nand NAND2_1697 (N6656, N1482, N6118);
  nand NAND2_1698 (N6657, N1485, N6120);
  nand NAND2_1699 (N6658, N3789, N6121);
  nand NAND2_1700 (N6659, N5039, N6123);
  nand NAND2_1701 (N6660, N5036, N6124);
  nand NAND2_1702 (N6661, N3792, N6126);
  nand NAND2_1703 (N6668, N3816, N6135);
  nand NAND2_1704 (N6677, N5071, N6148);
  nand NAND2_1705 (N6678, N5068, N6149);
  nand NAND2_1706 (N6679, N5077, N6150);
  nand NAND2_1707 (N6680, N5074, N6151);
  nand NAND2_1708 (N6681, N5083, N6152);
  nand NAND2_1709 (N6682, N5080, N6153);
  nand NAND2_1710 (N6683, N5089, N6154);
  nand NAND2_1711 (N6684, N5086, N6155);
  nand NAND2_1712 (N6685, N3846, N6156);
  nand NAND2_1713 (N6686, N3849, N6158);
  nand NAND2_1714 (N6687, N3852, N6160);
  nand NAND2_1715 (N6688, N5104, N6162);
  nand NAND2_1716 (N6689, N5101, N6163);
  nand NAND2_1717 (N6690, N3855, N6165);
  nand NAND2_1718 (N6702, N5117, N6181);
  nand NAND2_1719 (N6703, N5114, N6182);
  nand NAND2_1720 (N6704, N5123, N6183);
  nand NAND2_1721 (N6705, N5120, N6184);
  nand NAND2_1722 (N6706, N3891, N6185);
  nand NAND2_1723 (N6707, N5144, N6187);
  nand NAND2_1724 (N6708, N5141, N6188);
  nand NAND2_1725 (N6709, N5150, N6189);
  nand NAND2_1726 (N6710, N5147, N6190);
  nand NAND2_1727 (N6711, N1708, N6191);
  nand NAND2_1728 (N6712, N2231, N6193);
  nand NAND2_1729 (N6729, N4961, N6223);
  nand NAND2_1730 (N6730, N4958, N6224);
  nand NAND2_1731 (N6731, N4967, N6225);
  nand NAND2_1732 (N6732, N4964, N6226);
  nand NAND2_1733 (N6733, N4988, N6227);
  nand NAND2_1734 (N6734, N4985, N6228);
  nand NAND2_1735 (N6735, N4994, N6229);
  nand NAND2_1736 (N6736, N4991, N6230);
  nand NAND2_1737 (N6741, N5055, N6239);
  nand NAND2_1738 (N6742, N5052, N6240);
  nand NAND2_1739 (N6743, N5061, N6241);
  nand NAND2_1740 (N6744, N5058, N6242);
  nand NAND2_1741 (N6751, N5129, N6255);
  nand NAND2_1742 (N6752, N5126, N6256);
  nand NAND2_1743 (N6753, N5135, N6257);
  nand NAND2_1744 (N6754, N5132, N6258);
  nand NAND2_1745 (N6755, N5156, N6259);
  nand NAND2_1746 (N6756, N5153, N6260);
  nand NAND2_1747 (N6757, N5162, N6261);
  nand NAND2_1748 (N6758, N5159, N6262);
  not NOT1_1749 (N6761, N5892);
  and AND5_1750 (N6762, N5683, N5670, N5654, N5640, N5632);
  and AND2_1751 (N6766, N5632, N3097);
  and AND3_1752 (N6767, N5640, N5632, N3101);
  and AND4_1753 (N6768, N5654, N5632, N3107, N5640);
  and AND5_1754 (N6769, N5670, N5654, N5632, N3114, N5640);
  and AND2_1755 (N6770, N5640, N3101);
  and AND3_1756 (N6771, N5654, N3107, N5640);
  and AND4_1757 (N6772, N5670, N5654, N3114, N5640);
  and AND4_1758 (N6773, N5683, N5654, N5640, N5670);
  and AND2_1759 (N6774, N5640, N3101);
  and AND3_1760 (N6775, N5654, N3107, N5640);
  and AND4_1761 (N6776, N5670, N5654, N3114, N5640);
  and AND2_1762 (N6777, N5654, N3107);
  and AND3_1763 (N6778, N5670, N5654, N3114);
  and AND3_1764 (N6779, N5683, N5654, N5670);
  and AND2_1765 (N6780, N5654, N3107);
  and AND3_1766 (N6781, N5670, N5654, N3114);
  and AND2_1767 (N6782, N5670, N3114);
  and AND2_1768 (N6783, N5683, N5670);
  and AND5_1769 (N6784, N5697, N5728, N5707, N5690, N5718);
  and AND2_1770 (N6787, N5690, N3137);
  and AND3_1771 (N6788, N5697, N5690, N3140);
  and AND4_1772 (N6789, N5707, N5690, N3144, N5697);
  and AND5_1773 (N6790, N5718, N5707, N5690, N3149, N5697);
  and AND2_1774 (N6791, N5697, N3140);
  and AND3_1775 (N6792, N5707, N3144, N5697);
  and AND4_1776 (N6793, N5718, N5707, N3149, N5697);
  and AND2_1777 (N6794, N3144, N5707);
  and AND3_1778 (N6795, N5718, N5707, N3149);
  and AND2_1779 (N6796, N5718, N3149);
  not NOT1_1780 (N6797, N5736);
  not NOT1_1781 (N6800, N5740);
  not NOT1_1782 (N6803, N5747);
  not NOT1_1783 (N6806, N5751);
  not NOT1_1784 (N6809, N5758);
  not NOT1_1785 (N6812, N5762);
  buf BUFF1_1786 (N6815, N5744);
  buf BUFF1_1787 (N6818, N5744);
  buf BUFF1_1788 (N6821, N5755);
  buf BUFF1_1789 (N6824, N5755);
  buf BUFF1_1790 (N6827, N5766);
  buf BUFF1_1791 (N6830, N5766);
  and AND4_1792 (N6833, N5850, N5789, N5778, N5771);
  and AND2_1793 (N6836, N5771, N3169);
  and AND3_1794 (N6837, N5778, N5771, N3173);
  and AND4_1795 (N6838, N5789, N5771, N3178, N5778);
  and AND2_1796 (N6839, N5778, N3173);
  and AND3_1797 (N6840, N5789, N3178, N5778);
  and AND3_1798 (N6841, N5850, N5789, N5778);
  and AND2_1799 (N6842, N5778, N3173);
  and AND3_1800 (N6843, N5789, N3178, N5778);
  and AND2_1801 (N6844, N5789, N3178);
  and AND5_1802 (N6845, N5856, N5837, N5821, N5807, N5799);
  and AND2_1803 (N6848, N5799, N3185);
  and AND3_1804 (N6849, N5807, N5799, N3189);
  and AND4_1805 (N6850, N5821, N5799, N3195, N5807);
  and AND5_1806 (N6851, N5837, N5821, N5799, N3202, N5807);
  and AND2_1807 (N6852, N5807, N3189);
  and AND3_1808 (N6853, N5821, N3195, N5807);
  and AND4_1809 (N6854, N5837, N5821, N3202, N5807);
  and AND4_1810 (N6855, N5856, N5821, N5807, N5837);
  and AND2_1811 (N6856, N5807, N3189);
  and AND3_1812 (N6857, N5821, N3195, N5807);
  and AND4_1813 (N6858, N5837, N5821, N3202, N5807);
  and AND2_1814 (N6859, N5821, N3195);
  and AND3_1815 (N6860, N5837, N5821, N3202);
  and AND3_1816 (N6861, N5856, N5821, N5837);
  and AND2_1817 (N6862, N5821, N3195);
  and AND3_1818 (N6863, N5837, N5821, N3202);
  and AND2_1819 (N6864, N5837, N3202);
  and AND2_1820 (N6865, N5850, N5789);
  and AND2_1821 (N6866, N5856, N5837);
  and AND4_1822 (N6867, N5870, N5892, N5881, N5863);
  and AND2_1823 (N6870, N5863, N3211);
  and AND3_1824 (N6871, N5870, N5863, N3215);
  and AND4_1825 (N6872, N5881, N5863, N3221, N5870);
  and AND2_1826 (N6873, N5870, N3215);
  and AND3_1827 (N6874, N5881, N3221, N5870);
  and AND3_1828 (N6875, N5892, N5881, N5870);
  and AND2_1829 (N6876, N5870, N3215);
  and AND3_1830 (N6877, N3221, N5881, N5870);
  and AND2_1831 (N6878, N5881, N3221);
  and AND2_1832 (N6879, N5892, N5881);
  and AND2_1833 (N6880, N5881, N3221);
  and AND5_1834 (N6881, N5905, N5936, N5915, N5898, N5926);
  and AND2_1835 (N6884, N5898, N3229);
  and AND3_1836 (N6885, N5905, N5898, N3232);
  and AND4_1837 (N6886, N5915, N5898, N3236, N5905);
  and AND5_1838 (N6887, N5926, N5915, N5898, N3241, N5905);
  and AND2_1839 (N6888, N5905, N3232);
  and AND3_1840 (N6889, N5915, N3236, N5905);
  and AND4_1841 (N6890, N5926, N5915, N3241, N5905);
  and AND2_1842 (N6891, N3236, N5915);
  and AND3_1843 (N6892, N5926, N5915, N3241);
  and AND2_1844 (N6893, N5926, N3241);
  nand NAND2_1845 (N6894, N5944, N6540);
  nand NAND2_1846 (N6901, N5946, N6541);
  nand NAND2_1847 (N6912, N5948, N6542);
  nand NAND2_1848 (N6923, N5950, N6543);
  nand NAND2_1849 (N6929, N5952, N6544);
  nand NAND2_1850 (N6936, N5954, N6545);
  nand NAND2_1851 (N6946, N5956, N6546);
  nand NAND2_1852 (N6957, N5958, N6547);
  nand NAND2_1853 (N6967, N6204, N4575);
  not NOT1_1854 (N6968, N6204);
  not NOT1_1855 (N6969, N6207);
  nand NAND2_1856 (N6970, N5967, N6555);
  nand NAND2_1857 (N6977, N5969, N6556);
  nand NAND2_1858 (N6988, N5971, N6557);
  nand NAND2_1859 (N6998, N5973, N6558);
  nand NAND2_1860 (N7006, N5975, N6559);
  nand NAND2_1861 (N7020, N5977, N6560);
  nand NAND2_1862 (N7036, N5979, N6561);
  nand NAND2_1863 (N7049, N5989, N6569);
  nand NAND2_1864 (N7055, N6210, N4610);
  not NOT1_1865 (N7056, N6210);
  and AND4_1866 (N7057, N6021, N6000, N5996, N5991);
  and AND2_1867 (N7060, N5991, N3362);
  and AND3_1868 (N7061, N5996, N5991, N3363);
  and AND4_1869 (N7062, N6000, N5991, N3364, N5996);
  and AND5_1870 (N7063, N6022, N6018, N6014, N6009, N6003);
  and AND2_1871 (N7064, N6003, N3366);
  and AND3_1872 (N7065, N6009, N6003, N3367);
  and AND4_1873 (N7066, N6014, N6003, N3368, N6009);
  and AND5_1874 (N7067, N6018, N6014, N6003, N3369, N6009);
  nand NAND2_1875 (N7068, N6594, N6024);
  nand NAND2_1876 (N7073, N6595, N6026);
  nand NAND2_1877 (N7077, N6596, N6028);
  nand NAND2_1878 (N7080, N6597, N6030);
  nand NAND2_1879 (N7086, N6598, N6599);
  nand NAND2_1880 (N7091, N6600, N6601);
  nand NAND2_1881 (N7095, N6602, N6603);
  nand NAND2_1882 (N7098, N6604, N6038);
  nand NAND2_1883 (N7099, N6605, N6606);
  and AND5_1884 (N7100, N6059, N6056, N6052, N6047, N6041);
  and AND2_1885 (N7103, N6041, N3371);
  and AND3_1886 (N7104, N6047, N6041, N3372);
  and AND4_1887 (N7105, N6052, N6041, N3373, N6047);
  and AND5_1888 (N7106, N6056, N6052, N6041, N3374, N6047);
  nand NAND2_1889 (N7107, N6060, N6621);
  nand NAND2_1890 (N7114, N6062, N6622);
  nand NAND2_1891 (N7125, N6064, N6623);
  nand NAND2_1892 (N7136, N6066, N6624);
  nand NAND2_1893 (N7142, N6068, N6625);
  nand NAND2_1894 (N7149, N6070, N6626);
  nand NAND2_1895 (N7159, N6072, N6627);
  nand NAND2_1896 (N7170, N6074, N6628);
  nand NAND2_1897 (N7180, N6076, N6629);
  not NOT1_1898 (N7187, N6220);
  not NOT1_1899 (N7188, N6079);
  not NOT1_1900 (N7191, N6083);
  nand NAND2_1901 (N7194, N6639, N6091);
  nand NAND2_1902 (N7198, N6640, N6641);
  nand NAND2_1903 (N7202, N6642, N6643);
  nand NAND2_1904 (N7205, N6644, N6097);
  nand NAND2_1905 (N7209, N6645, N6646);
  nand NAND2_1906 (N7213, N6647, N6648);
  buf BUFF1_1907 (N7216, N6087);
  buf BUFF1_1908 (N7219, N6087);
  nand NAND2_1909 (N7222, N6103, N6649);
  nand NAND2_1910 (N7229, N6105, N6650);
  nand NAND2_1911 (N7240, N6107, N6651);
  nand NAND2_1912 (N7250, N6109, N6652);
  nand NAND2_1913 (N7258, N6111, N6653);
  nand NAND2_1914 (N7272, N6113, N6654);
  nand NAND2_1915 (N7288, N6115, N6655);
  nand NAND2_1916 (N7301, N6117, N6656);
  nand NAND2_1917 (N7307, N6119, N6657);
  nand NAND2_1918 (N7314, N6658, N6122);
  nand NAND2_1919 (N7318, N6659, N6660);
  nand NAND2_1920 (N7322, N6125, N6661);
  not NOT1_1921 (N7325, N6127);
  not NOT1_1922 (N7328, N6131);
  nand NAND2_1923 (N7331, N6668, N6136);
  not NOT1_1924 (N7334, N6137);
  not NOT1_1925 (N7337, N6141);
  buf BUFF1_1926 (N7340, N6145);
  buf BUFF1_1927 (N7343, N6145);
  nand NAND2_1928 (N7346, N6677, N6678);
  nand NAND2_1929 (N7351, N6679, N6680);
  nand NAND2_1930 (N7355, N6681, N6682);
  nand NAND2_1931 (N7358, N6683, N6684);
  nand NAND2_1932 (N7364, N6685, N6157);
  nand NAND2_1933 (N7369, N6686, N6159);
  nand NAND2_1934 (N7373, N6687, N6161);
  nand NAND2_1935 (N7376, N6688, N6689);
  nand NAND2_1936 (N7377, N6164, N6690);
  not NOT1_1937 (N7378, N6166);
  not NOT1_1938 (N7381, N6170);
  not NOT1_1939 (N7384, N6177);
  nand NAND2_1940 (N7387, N6702, N6703);
  nand NAND2_1941 (N7391, N6704, N6705);
  nand NAND2_1942 (N7394, N6706, N6186);
  nand NAND2_1943 (N7398, N6707, N6708);
  nand NAND2_1944 (N7402, N6709, N6710);
  buf BUFF1_1945 (N7405, N6174);
  buf BUFF1_1946 (N7408, N6174);
  buf BUFF1_1947 (N7411, N5936);
  buf BUFF1_1948 (N7414, N5898);
  buf BUFF1_1949 (N7417, N5905);
  buf BUFF1_1950 (N7420, N5915);
  buf BUFF1_1951 (N7423, N5926);
  buf BUFF1_1952 (N7426, N5728);
  buf BUFF1_1953 (N7429, N5690);
  buf BUFF1_1954 (N7432, N5697);
  buf BUFF1_1955 (N7435, N5707);
  buf BUFF1_1956 (N7438, N5718);
  nand NAND2_1957 (N7441, N6192, N6711);
  nand NAND2_1958 (N7444, N6194, N6712);
  buf BUFF1_1959 (N7447, N5683);
  buf BUFF1_1960 (N7450, N5670);
  buf BUFF1_1961 (N7453, N5632);
  buf BUFF1_1962 (N7456, N5654);
  buf BUFF1_1963 (N7459, N5640);
  buf BUFF1_1964 (N7462, N5640);
  buf BUFF1_1965 (N7465, N5683);
  buf BUFF1_1966 (N7468, N5670);
  buf BUFF1_1967 (N7471, N5632);
  buf BUFF1_1968 (N7474, N5654);
  not NOT1_1969 (N7477, N6196);
  not NOT1_1970 (N7478, N6199);
  buf BUFF1_1971 (N7479, N5850);
  buf BUFF1_1972 (N7482, N5789);
  buf BUFF1_1973 (N7485, N5771);
  buf BUFF1_1974 (N7488, N5778);
  buf BUFF1_1975 (N7491, N5850);
  buf BUFF1_1976 (N7494, N5789);
  buf BUFF1_1977 (N7497, N5771);
  buf BUFF1_1978 (N7500, N5778);
  buf BUFF1_1979 (N7503, N5856);
  buf BUFF1_1980 (N7506, N5837);
  buf BUFF1_1981 (N7509, N5799);
  buf BUFF1_1982 (N7512, N5821);
  buf BUFF1_1983 (N7515, N5807);
  buf BUFF1_1984 (N7518, N5807);
  buf BUFF1_1985 (N7521, N5856);
  buf BUFF1_1986 (N7524, N5837);
  buf BUFF1_1987 (N7527, N5799);
  buf BUFF1_1988 (N7530, N5821);
  buf BUFF1_1989 (N7533, N5863);
  buf BUFF1_1990 (N7536, N5863);
  buf BUFF1_1991 (N7539, N5870);
  buf BUFF1_1992 (N7542, N5870);
  buf BUFF1_1993 (N7545, N5881);
  buf BUFF1_1994 (N7548, N5881);
  not NOT1_1995 (N7551, N6214);
  not NOT1_1996 (N7552, N6217);
  buf BUFF1_1997 (N7553, N5981);
  not NOT1_1998 (N7556, N6249);
  not NOT1_1999 (N7557, N6252);
  not NOT1_2000 (N7558, N6243);
  not NOT1_2001 (N7559, N6246);
  nand NAND2_2002 (N7560, N6731, N6732);
  nand NAND2_2003 (N7563, N6729, N6730);
  nand NAND2_2004 (N7566, N6735, N6736);
  nand NAND2_2005 (N7569, N6733, N6734);
  not NOT1_2006 (N7572, N6232);
  not NOT1_2007 (N7573, N6236);
  nand NAND2_2008 (N7574, N6743, N6744);
  nand NAND2_2009 (N7577, N6741, N6742);
  not NOT1_2010 (N7580, N6263);
  not NOT1_2011 (N7581, N6266);
  nand NAND2_2012 (N7582, N6753, N6754);
  nand NAND2_2013 (N7585, N6751, N6752);
  nand NAND2_2014 (N7588, N6757, N6758);
  nand NAND2_2015 (N7591, N6755, N6756);
  or OR5_2016 (N7609, N3096, N6766, N6767, N6768, N6769);
  or OR2_2017 (N7613, N3107, N6782);
  or OR5_2018 (N7620, N3136, N6787, N6788, N6789, N6790);
  or OR4_2019 (N7649, N3168, N6836, N6837, N6838);
  or OR2_2020 (N7650, N3173, N6844);
  or OR5_2021 (N7655, N3184, N6848, N6849, N6850, N6851);
  or OR2_2022 (N7659, N3195, N6864);
  or OR4_2023 (N7668, N3210, N6870, N6871, N6872);
  or OR5_2024 (N7671, N3228, N6884, N6885, N6886, N6887);
  nand NAND2_2025 (N7744, N3661, N6968);
  nand NAND2_2026 (N7822, N3664, N7056);
  or OR4_2027 (N7825, N3361, N7060, N7061, N7062);
  or OR5_2028 (N7826, N3365, N7064, N7065, N7066, N7067);
  or OR5_2029 (N7852, N3370, N7103, N7104, N7105, N7106);
  or OR4_2030 (N8114, N3101, N6777, N6778, N6779);
  or OR5_2031 (N8117, N3097, N6770, N6771, N6772, N6773);
  nor NOR3_2032 (N8131, N3101, N6780, N6781);
  nor NOR4_2033 (N8134, N3097, N6774, N6775, N6776);
  nand NAND2_2034 (N8144, N6199, N7477);
  nand NAND2_2035 (N8145, N6196, N7478);
  or OR4_2036 (N8146, N3169, N6839, N6840, N6841);
  nor NOR3_2037 (N8156, N3169, N6842, N6843);
  or OR4_2038 (N8166, N3189, N6859, N6860, N6861);
  or OR5_2039 (N8169, N3185, N6852, N6853, N6854, N6855);
  nor NOR3_2040 (N8183, N3189, N6862, N6863);
  nor NOR4_2041 (N8186, N3185, N6856, N6857, N6858);
  or OR4_2042 (N8196, N3211, N6873, N6874, N6875);
  nor NOR3_2043 (N8200, N3211, N6876, N6877);
  or OR3_2044 (N8204, N3215, N6878, N6879);
  nor NOR2_2045 (N8208, N3215, N6880);
  nand NAND2_2046 (N8216, N6252, N7556);
  nand NAND2_2047 (N8217, N6249, N7557);
  nand NAND2_2048 (N8218, N6246, N7558);
  nand NAND2_2049 (N8219, N6243, N7559);
  nand NAND2_2050 (N8232, N6266, N7580);
  nand NAND2_2051 (N8233, N6263, N7581);
  not NOT1_2052 (N8242, N7411);
  not NOT1_2053 (N8243, N7414);
  not NOT1_2054 (N8244, N7417);
  not NOT1_2055 (N8245, N7420);
  not NOT1_2056 (N8246, N7423);
  not NOT1_2057 (N8247, N7426);
  not NOT1_2058 (N8248, N7429);
  not NOT1_2059 (N8249, N7432);
  not NOT1_2060 (N8250, N7435);
  not NOT1_2061 (N8251, N7438);
  not NOT1_2062 (N8252, N7136);
  not NOT1_2063 (N8253, N6923);
  not NOT1_2064 (N8254, N6762);
  not NOT1_2065 (N8260, N7459);
  not NOT1_2066 (N8261, N7462);
  and AND2_2067 (N8262, N3122, N6762);
  and AND2_2068 (N8269, N3155, N6784);
  not NOT1_2069 (N8274, N6815);
  not NOT1_2070 (N8275, N6818);
  not NOT1_2071 (N8276, N6821);
  not NOT1_2072 (N8277, N6824);
  not NOT1_2073 (N8278, N6827);
  not NOT1_2074 (N8279, N6830);
  and AND3_2075 (N8280, N5740, N5736, N6815);
  and AND3_2076 (N8281, N6800, N6797, N6818);
  and AND3_2077 (N8282, N5751, N5747, N6821);
  and AND3_2078 (N8283, N6806, N6803, N6824);
  and AND3_2079 (N8284, N5762, N5758, N6827);
  and AND3_2080 (N8285, N6812, N6809, N6830);
  not NOT1_2081 (N8288, N6845);
  not NOT1_2082 (N8294, N7488);
  not NOT1_2083 (N8295, N7500);
  not NOT1_2084 (N8296, N7515);
  not NOT1_2085 (N8297, N7518);
  and AND2_2086 (N8298, N6833, N6845);
  and AND2_2087 (N8307, N6867, N6881);
  not NOT1_2088 (N8315, N7533);
  not NOT1_2089 (N8317, N7536);
  not NOT1_2090 (N8319, N7539);
  not NOT1_2091 (N8321, N7542);
  nand NAND2_2092 (N8322, N7545, N4543);
  not NOT1_2093 (N8323, N7545);
  nand NAND2_2094 (N8324, N7548, N5943);
  not NOT1_2095 (N8325, N7548);
  nand NAND2_2096 (N8326, N6967, N7744);
  and AND4_2097 (N8333, N6901, N6923, N6912, N6894);
  and AND2_2098 (N8337, N6894, N4545);
  and AND3_2099 (N8338, N6901, N6894, N4549);
  and AND4_2100 (N8339, N6912, N6894, N4555, N6901);
  and AND2_2101 (N8340, N6901, N4549);
  and AND3_2102 (N8341, N6912, N4555, N6901);
  and AND3_2103 (N8342, N6923, N6912, N6901);
  and AND2_2104 (N8343, N6901, N4549);
  and AND3_2105 (N8344, N4555, N6912, N6901);
  and AND2_2106 (N8345, N6912, N4555);
  and AND2_2107 (N8346, N6923, N6912);
  and AND2_2108 (N8347, N6912, N4555);
  and AND2_2109 (N8348, N6929, N4563);
  and AND3_2110 (N8349, N6936, N6929, N4566);
  and AND4_2111 (N8350, N6946, N6929, N4570, N6936);
  and AND5_2112 (N8351, N6957, N6946, N6929, N5960, N6936);
  and AND2_2113 (N8352, N6936, N4566);
  and AND3_2114 (N8353, N6946, N4570, N6936);
  and AND4_2115 (N8354, N6957, N6946, N5960, N6936);
  and AND2_2116 (N8355, N4570, N6946);
  and AND3_2117 (N8356, N6957, N6946, N5960);
  and AND2_2118 (N8357, N6957, N5960);
  nand NAND2_2119 (N8358, N7055, N7822);
  and AND4_2120 (N8365, N7049, N6988, N6977, N6970);
  and AND2_2121 (N8369, N6970, N4577);
  and AND3_2122 (N8370, N6977, N6970, N4581);
  and AND4_2123 (N8371, N6988, N6970, N4586, N6977);
  and AND2_2124 (N8372, N6977, N4581);
  and AND3_2125 (N8373, N6988, N4586, N6977);
  and AND3_2126 (N8374, N7049, N6988, N6977);
  and AND2_2127 (N8375, N6977, N4581);
  and AND3_2128 (N8376, N6988, N4586, N6977);
  and AND2_2129 (N8377, N6988, N4586);
  and AND2_2130 (N8378, N6998, N4593);
  and AND3_2131 (N8379, N7006, N6998, N4597);
  and AND4_2132 (N8380, N7020, N6998, N4603, N7006);
  and AND5_2133 (N8381, N7036, N7020, N6998, N5981, N7006);
  and AND2_2134 (N8382, N7006, N4597);
  and AND3_2135 (N8383, N7020, N4603, N7006);
  and AND4_2136 (N8384, N7036, N7020, N5981, N7006);
  and AND2_2137 (N8385, N7006, N4597);
  and AND3_2138 (N8386, N7020, N4603, N7006);
  and AND4_2139 (N8387, N7036, N7020, N5981, N7006);
  and AND2_2140 (N8388, N7020, N4603);
  and AND3_2141 (N8389, N7036, N7020, N5981);
  and AND2_2142 (N8390, N7020, N4603);
  and AND3_2143 (N8391, N7036, N7020, N5981);
  and AND2_2144 (N8392, N7036, N5981);
  and AND2_2145 (N8393, N7049, N6988);
  and AND2_2146 (N8394, N7057, N7063);
  and AND2_2147 (N8404, N7057, N7826);
  and AND4_2148 (N8405, N7098, N7077, N7073, N7068);
  and AND2_2149 (N8409, N7068, N4632);
  and AND3_2150 (N8410, N7073, N7068, N4634);
  and AND4_2151 (N8411, N7077, N7068, N4635, N7073);
  and AND5_2152 (N8412, N7099, N7095, N7091, N7086, N7080);
  and AND2_2153 (N8415, N7080, N4638);
  and AND3_2154 (N8416, N7086, N7080, N4639);
  and AND4_2155 (N8417, N7091, N7080, N4640, N7086);
  and AND5_2156 (N8418, N7095, N7091, N7080, N4641, N7086);
  and AND2_2157 (N8421, N3375, N7100);
  and AND4_2158 (N8430, N7114, N7136, N7125, N7107);
  and AND2_2159 (N8433, N7107, N4657);
  and AND3_2160 (N8434, N7114, N7107, N4661);
  and AND4_2161 (N8435, N7125, N7107, N4667, N7114);
  and AND2_2162 (N8436, N7114, N4661);
  and AND3_2163 (N8437, N7125, N4667, N7114);
  and AND3_2164 (N8438, N7136, N7125, N7114);
  and AND2_2165 (N8439, N7114, N4661);
  and AND3_2166 (N8440, N4667, N7125, N7114);
  and AND2_2167 (N8441, N7125, N4667);
  and AND2_2168 (N8442, N7136, N7125);
  and AND2_2169 (N8443, N7125, N4667);
  and AND5_2170 (N8444, N7149, N7180, N7159, N7142, N7170);
  and AND2_2171 (N8447, N7142, N4675);
  and AND3_2172 (N8448, N7149, N7142, N4678);
  and AND4_2173 (N8449, N7159, N7142, N4682, N7149);
  and AND5_2174 (N8450, N7170, N7159, N7142, N4687, N7149);
  and AND2_2175 (N8451, N7149, N4678);
  and AND3_2176 (N8452, N7159, N4682, N7149);
  and AND4_2177 (N8453, N7170, N7159, N4687, N7149);
  and AND2_2178 (N8454, N4682, N7159);
  and AND3_2179 (N8455, N7170, N7159, N4687);
  and AND2_2180 (N8456, N7170, N4687);
  not NOT1_2181 (N8457, N7194);
  not NOT1_2182 (N8460, N7198);
  not NOT1_2183 (N8463, N7205);
  not NOT1_2184 (N8466, N7209);
  not NOT1_2185 (N8469, N7216);
  not NOT1_2186 (N8470, N7219);
  buf BUFF1_2187 (N8471, N7202);
  buf BUFF1_2188 (N8474, N7202);
  buf BUFF1_2189 (N8477, N7213);
  buf BUFF1_2190 (N8480, N7213);
  and AND3_2191 (N8483, N6083, N6079, N7216);
  and AND3_2192 (N8484, N7191, N7188, N7219);
  and AND4_2193 (N8485, N7301, N7240, N7229, N7222);
  and AND2_2194 (N8488, N7222, N4702);
  and AND3_2195 (N8489, N7229, N7222, N4706);
  and AND4_2196 (N8490, N7240, N7222, N4711, N7229);
  and AND2_2197 (N8491, N7229, N4706);
  and AND3_2198 (N8492, N7240, N4711, N7229);
  and AND3_2199 (N8493, N7301, N7240, N7229);
  and AND2_2200 (N8494, N7229, N4706);
  and AND3_2201 (N8495, N7240, N4711, N7229);
  and AND2_2202 (N8496, N7240, N4711);
  and AND5_2203 (N8497, N7307, N7288, N7272, N7258, N7250);
  and AND2_2204 (N8500, N7250, N4718);
  and AND3_2205 (N8501, N7258, N7250, N4722);
  and AND4_2206 (N8502, N7272, N7250, N4728, N7258);
  and AND5_2207 (N8503, N7288, N7272, N7250, N4735, N7258);
  and AND2_2208 (N8504, N7258, N4722);
  and AND3_2209 (N8505, N7272, N4728, N7258);
  and AND4_2210 (N8506, N7288, N7272, N4735, N7258);
  and AND4_2211 (N8507, N7307, N7272, N7258, N7288);
  and AND2_2212 (N8508, N7258, N4722);
  and AND3_2213 (N8509, N7272, N4728, N7258);
  and AND4_2214 (N8510, N7288, N7272, N4735, N7258);
  and AND2_2215 (N8511, N7272, N4728);
  and AND3_2216 (N8512, N7288, N7272, N4735);
  and AND3_2217 (N8513, N7307, N7272, N7288);
  and AND2_2218 (N8514, N7272, N4728);
  and AND3_2219 (N8515, N7288, N7272, N4735);
  and AND2_2220 (N8516, N7288, N4735);
  and AND2_2221 (N8517, N7301, N7240);
  and AND2_2222 (N8518, N7307, N7288);
  not NOT1_2223 (N8519, N7314);
  not NOT1_2224 (N8522, N7318);
  buf BUFF1_2225 (N8525, N7322);
  buf BUFF1_2226 (N8528, N7322);
  buf BUFF1_2227 (N8531, N7331);
  buf BUFF1_2228 (N8534, N7331);
  not NOT1_2229 (N8537, N7340);
  not NOT1_2230 (N8538, N7343);
  and AND3_2231 (N8539, N6141, N6137, N7340);
  and AND3_2232 (N8540, N7337, N7334, N7343);
  and AND4_2233 (N8541, N7376, N7355, N7351, N7346);
  and AND2_2234 (N8545, N7346, N4757);
  and AND3_2235 (N8546, N7351, N7346, N4758);
  and AND4_2236 (N8547, N7355, N7346, N4759, N7351);
  and AND5_2237 (N8548, N7377, N7373, N7369, N7364, N7358);
  and AND2_2238 (N8551, N7358, N4762);
  and AND3_2239 (N8552, N7364, N7358, N4764);
  and AND4_2240 (N8553, N7369, N7358, N4766, N7364);
  and AND5_2241 (N8554, N7373, N7369, N7358, N4767, N7364);
  not NOT1_2242 (N8555, N7387);
  not NOT1_2243 (N8558, N7394);
  not NOT1_2244 (N8561, N7398);
  not NOT1_2245 (N8564, N7405);
  not NOT1_2246 (N8565, N7408);
  buf BUFF1_2247 (N8566, N7391);
  buf BUFF1_2248 (N8569, N7391);
  buf BUFF1_2249 (N8572, N7402);
  buf BUFF1_2250 (N8575, N7402);
  and AND3_2251 (N8578, N6170, N6166, N7405);
  and AND3_2252 (N8579, N7381, N7378, N7408);
  buf BUFF1_2253 (N8580, N7180);
  buf BUFF1_2254 (N8583, N7142);
  buf BUFF1_2255 (N8586, N7149);
  buf BUFF1_2256 (N8589, N7159);
  buf BUFF1_2257 (N8592, N7170);
  buf BUFF1_2258 (N8595, N6929);
  buf BUFF1_2259 (N8598, N6936);
  buf BUFF1_2260 (N8601, N6946);
  buf BUFF1_2261 (N8604, N6957);
  not NOT1_2262 (N8607, N7441);
  nand NAND2_2263 (N8608, N7441, N5469);
  not NOT1_2264 (N8609, N7444);
  nand NAND2_2265 (N8610, N7444, N4793);
  not NOT1_2266 (N8615, N7447);
  not NOT1_2267 (N8616, N7450);
  not NOT1_2268 (N8617, N7453);
  not NOT1_2269 (N8618, N7456);
  not NOT1_2270 (N8619, N7474);
  not NOT1_2271 (N8624, N7465);
  not NOT1_2272 (N8625, N7468);
  not NOT1_2273 (N8626, N7471);
  nand NAND2_2274 (N8627, N8144, N8145);
  not NOT1_2275 (N8632, N7479);
  not NOT1_2276 (N8633, N7482);
  not NOT1_2277 (N8634, N7485);
  not NOT1_2278 (N8637, N7491);
  not NOT1_2279 (N8638, N7494);
  not NOT1_2280 (N8639, N7497);
  not NOT1_2281 (N8644, N7503);
  not NOT1_2282 (N8645, N7506);
  not NOT1_2283 (N8646, N7509);
  not NOT1_2284 (N8647, N7512);
  not NOT1_2285 (N8648, N7530);
  not NOT1_2286 (N8653, N7521);
  not NOT1_2287 (N8654, N7524);
  not NOT1_2288 (N8655, N7527);
  buf BUFF1_2289 (N8660, N6894);
  buf BUFF1_2290 (N8663, N6894);
  buf BUFF1_2291 (N8666, N6901);
  buf BUFF1_2292 (N8669, N6901);
  buf BUFF1_2293 (N8672, N6912);
  buf BUFF1_2294 (N8675, N6912);
  buf BUFF1_2295 (N8678, N7049);
  buf BUFF1_2296 (N8681, N6988);
  buf BUFF1_2297 (N8684, N6970);
  buf BUFF1_2298 (N8687, N6977);
  buf BUFF1_2299 (N8690, N7049);
  buf BUFF1_2300 (N8693, N6988);
  buf BUFF1_2301 (N8696, N6970);
  buf BUFF1_2302 (N8699, N6977);
  buf BUFF1_2303 (N8702, N7036);
  buf BUFF1_2304 (N8705, N6998);
  buf BUFF1_2305 (N8708, N7020);
  buf BUFF1_2306 (N8711, N7006);
  buf BUFF1_2307 (N8714, N7006);
  not NOT1_2308 (N8717, N7553);
  buf BUFF1_2309 (N8718, N7036);
  buf BUFF1_2310 (N8721, N6998);
  buf BUFF1_2311 (N8724, N7020);
  nand NAND2_2312 (N8727, N8216, N8217);
  nand NAND2_2313 (N8730, N8218, N8219);
  not NOT1_2314 (N8733, N7574);
  not NOT1_2315 (N8734, N7577);
  buf BUFF1_2316 (N8735, N7107);
  buf BUFF1_2317 (N8738, N7107);
  buf BUFF1_2318 (N8741, N7114);
  buf BUFF1_2319 (N8744, N7114);
  buf BUFF1_2320 (N8747, N7125);
  buf BUFF1_2321 (N8750, N7125);
  not NOT1_2322 (N8753, N7560);
  not NOT1_2323 (N8754, N7563);
  not NOT1_2324 (N8755, N7566);
  not NOT1_2325 (N8756, N7569);
  buf BUFF1_2326 (N8757, N7301);
  buf BUFF1_2327 (N8760, N7240);
  buf BUFF1_2328 (N8763, N7222);
  buf BUFF1_2329 (N8766, N7229);
  buf BUFF1_2330 (N8769, N7301);
  buf BUFF1_2331 (N8772, N7240);
  buf BUFF1_2332 (N8775, N7222);
  buf BUFF1_2333 (N8778, N7229);
  buf BUFF1_2334 (N8781, N7307);
  buf BUFF1_2335 (N8784, N7288);
  buf BUFF1_2336 (N8787, N7250);
  buf BUFF1_2337 (N8790, N7272);
  buf BUFF1_2338 (N8793, N7258);
  buf BUFF1_2339 (N8796, N7258);
  buf BUFF1_2340 (N8799, N7307);
  buf BUFF1_2341 (N8802, N7288);
  buf BUFF1_2342 (N8805, N7250);
  buf BUFF1_2343 (N8808, N7272);
  nand NAND2_2344 (N8811, N8232, N8233);
  not NOT1_2345 (N8814, N7588);
  not NOT1_2346 (N8815, N7591);
  not NOT1_2347 (N8816, N7582);
  not NOT1_2348 (N8817, N7585);
  and AND2_2349 (N8818, N7620, N3155);
  and AND2_2350 (N8840, N3122, N7609);
  not NOT1_2351 (N8857, N7609);
  and AND3_2352 (N8861, N6797, N5740, N8274);
  and AND3_2353 (N8862, N5736, N6800, N8275);
  and AND3_2354 (N8863, N6803, N5751, N8276);
  and AND3_2355 (N8864, N5747, N6806, N8277);
  and AND3_2356 (N8865, N6809, N5762, N8278);
  and AND3_2357 (N8866, N5758, N6812, N8279);
  not NOT1_2358 (N8871, N7655);
  and AND2_2359 (N8874, N6833, N7655);
  and AND2_2360 (N8878, N7671, N6867);
  not NOT1_2361 (N8879, N8196);
  nand NAND2_2362 (N8880, N8196, N8315);
  not NOT1_2363 (N8881, N8200);
  nand NAND2_2364 (N8882, N8200, N8317);
  not NOT1_2365 (N8883, N8204);
  nand NAND2_2366 (N8884, N8204, N8319);
  not NOT1_2367 (N8885, N8208);
  nand NAND2_2368 (N8886, N8208, N8321);
  nand NAND2_2369 (N8887, N3658, N8323);
  nand NAND2_2370 (N8888, N4817, N8325);
  or OR4_2371 (N8898, N4544, N8337, N8338, N8339);
  or OR5_2372 (N8902, N4562, N8348, N8349, N8350, N8351);
  or OR4_2373 (N8920, N4576, N8369, N8370, N8371);
  or OR2_2374 (N8924, N4581, N8377);
  or OR5_2375 (N8927, N4592, N8378, N8379, N8380, N8381);
  or OR2_2376 (N8931, N4603, N8392);
  or OR2_2377 (N8943, N7825, N8404);
  or OR4_2378 (N8950, N4630, N8409, N8410, N8411);
  or OR5_2379 (N8956, N4637, N8415, N8416, N8417, N8418);
  not NOT1_2380 (N8959, N7852);
  and AND2_2381 (N8960, N3375, N7852);
  or OR4_2382 (N8963, N4656, N8433, N8434, N8435);
  or OR5_2383 (N8966, N4674, N8447, N8448, N8449, N8450);
  and AND3_2384 (N8991, N7188, N6083, N8469);
  and AND3_2385 (N8992, N6079, N7191, N8470);
  or OR4_2386 (N8995, N4701, N8488, N8489, N8490);
  or OR2_2387 (N8996, N4706, N8496);
  or OR5_2388 (N9001, N4717, N8500, N8501, N8502, N8503);
  or OR2_2389 (N9005, N4728, N8516);
  and AND3_2390 (N9024, N7334, N6141, N8537);
  and AND3_2391 (N9025, N6137, N7337, N8538);
  or OR4_2392 (N9029, N4756, N8545, N8546, N8547);
  or OR5_2393 (N9035, N4760, N8551, N8552, N8553, N8554);
  and AND3_2394 (N9053, N7378, N6170, N8564);
  and AND3_2395 (N9054, N6166, N7381, N8565);
  nand NAND2_2396 (N9064, N4303, N8607);
  nand NAND2_2397 (N9065, N3507, N8609);
  not NOT1_2398 (N9066, N8114);
  nand NAND2_2399 (N9067, N8114, N4795);
  or OR2_2400 (N9068, N7613, N6783);
  not NOT1_2401 (N9071, N8117);
  not NOT1_2402 (N9072, N8131);
  nand NAND2_2403 (N9073, N8131, N6195);
  not NOT1_2404 (N9074, N7613);
  not NOT1_2405 (N9077, N8134);
  or OR2_2406 (N9079, N7650, N6865);
  not NOT1_2407 (N9082, N8146);
  not NOT1_2408 (N9083, N7650);
  not NOT1_2409 (N9086, N8156);
  not NOT1_2410 (N9087, N8166);
  nand NAND2_2411 (N9088, N8166, N4813);
  or OR2_2412 (N9089, N7659, N6866);
  not NOT1_2413 (N9092, N8169);
  not NOT1_2414 (N9093, N8183);
  nand NAND2_2415 (N9094, N8183, N6203);
  not NOT1_2416 (N9095, N7659);
  not NOT1_2417 (N9098, N8186);
  or OR4_2418 (N9099, N4545, N8340, N8341, N8342);
  nor NOR3_2419 (N9103, N4545, N8343, N8344);
  or OR3_2420 (N9107, N4549, N8345, N8346);
  nor NOR2_2421 (N9111, N4549, N8347);
  or OR4_2422 (N9117, N4577, N8372, N8373, N8374);
  nor NOR3_2423 (N9127, N4577, N8375, N8376);
  nor NOR3_2424 (N9146, N4597, N8390, N8391);
  nor NOR4_2425 (N9149, N4593, N8385, N8386, N8387);
  nand NAND2_2426 (N9159, N7577, N8733);
  nand NAND2_2427 (N9160, N7574, N8734);
  or OR4_2428 (N9161, N4657, N8436, N8437, N8438);
  nor NOR3_2429 (N9165, N4657, N8439, N8440);
  or OR3_2430 (N9169, N4661, N8441, N8442);
  nor NOR2_2431 (N9173, N4661, N8443);
  nand NAND2_2432 (N9179, N7563, N8753);
  nand NAND2_2433 (N9180, N7560, N8754);
  nand NAND2_2434 (N9181, N7569, N8755);
  nand NAND2_2435 (N9182, N7566, N8756);
  or OR4_2436 (N9183, N4702, N8491, N8492, N8493);
  nor NOR3_2437 (N9193, N4702, N8494, N8495);
  or OR4_2438 (N9203, N4722, N8511, N8512, N8513);
  or OR5_2439 (N9206, N4718, N8504, N8505, N8506, N8507);
  nor NOR3_2440 (N9220, N4722, N8514, N8515);
  nor NOR4_2441 (N9223, N4718, N8508, N8509, N8510);
  nand NAND2_2442 (N9234, N7591, N8814);
  nand NAND2_2443 (N9235, N7588, N8815);
  nand NAND2_2444 (N9236, N7585, N8816);
  nand NAND2_2445 (N9237, N7582, N8817);
  or OR2_2446 (N9238, N3159, N8818);
  or OR2_2447 (N9242, N3126, N8840);
  nand NAND2_2448 (N9243, N8324, N8888);
  not NOT1_2449 (N9244, N8580);
  not NOT1_2450 (N9245, N8583);
  not NOT1_2451 (N9246, N8586);
  not NOT1_2452 (N9247, N8589);
  not NOT1_2453 (N9248, N8592);
  not NOT1_2454 (N9249, N8595);
  not NOT1_2455 (N9250, N8598);
  not NOT1_2456 (N9251, N8601);
  not NOT1_2457 (N9252, N8604);
  nor NOR2_2458 (N9256, N8861, N8280);
  nor NOR2_2459 (N9257, N8862, N8281);
  nor NOR2_2460 (N9258, N8863, N8282);
  nor NOR2_2461 (N9259, N8864, N8283);
  nor NOR2_2462 (N9260, N8865, N8284);
  nor NOR2_2463 (N9261, N8866, N8285);
  not NOT1_2464 (N9262, N8627);
  or OR2_2465 (N9265, N7649, N8874);
  or OR2_2466 (N9268, N7668, N8878);
  nand NAND2_2467 (N9271, N7533, N8879);
  nand NAND2_2468 (N9272, N7536, N8881);
  nand NAND2_2469 (N9273, N7539, N8883);
  nand NAND2_2470 (N9274, N7542, N8885);
  nand NAND2_2471 (N9275, N8322, N8887);
  not NOT1_2472 (N9276, N8333);
  and AND5_2473 (N9280, N6936, N8326, N6946, N6929, N6957);
  and AND5_2474 (N9285, N367, N8326, N6946, N6957, N6936);
  and AND4_2475 (N9286, N367, N8326, N6946, N6957);
  and AND3_2476 (N9287, N367, N8326, N6957);
  and AND2_2477 (N9288, N367, N8326);
  not NOT1_2478 (N9290, N8660);
  not NOT1_2479 (N9292, N8663);
  not NOT1_2480 (N9294, N8666);
  not NOT1_2481 (N9296, N8669);
  nand NAND2_2482 (N9297, N8672, N5966);
  not NOT1_2483 (N9298, N8672);
  nand NAND2_2484 (N9299, N8675, N6969);
  not NOT1_2485 (N9300, N8675);
  not NOT1_2486 (N9301, N8365);
  and AND5_2487 (N9307, N8358, N7036, N7020, N7006, N6998);
  and AND4_2488 (N9314, N8358, N7020, N7006, N7036);
  and AND3_2489 (N9315, N8358, N7020, N7036);
  and AND2_2490 (N9318, N8358, N7036);
  not NOT1_2491 (N9319, N8687);
  not NOT1_2492 (N9320, N8699);
  not NOT1_2493 (N9321, N8711);
  not NOT1_2494 (N9322, N8714);
  not NOT1_2495 (N9323, N8727);
  not NOT1_2496 (N9324, N8730);
  not NOT1_2497 (N9326, N8405);
  and AND2_2498 (N9332, N8405, N8412);
  or OR2_2499 (N9339, N4193, N8960);
  and AND2_2500 (N9344, N8430, N8444);
  not NOT1_2501 (N9352, N8735);
  not NOT1_2502 (N9354, N8738);
  not NOT1_2503 (N9356, N8741);
  not NOT1_2504 (N9358, N8744);
  nand NAND2_2505 (N9359, N8747, N6078);
  not NOT1_2506 (N9360, N8747);
  nand NAND2_2507 (N9361, N8750, N7187);
  not NOT1_2508 (N9362, N8750);
  not NOT1_2509 (N9363, N8471);
  not NOT1_2510 (N9364, N8474);
  not NOT1_2511 (N9365, N8477);
  not NOT1_2512 (N9366, N8480);
  nor NOR2_2513 (N9367, N8991, N8483);
  nor NOR2_2514 (N9368, N8992, N8484);
  and AND3_2515 (N9369, N7198, N7194, N8471);
  and AND3_2516 (N9370, N8460, N8457, N8474);
  and AND3_2517 (N9371, N7209, N7205, N8477);
  and AND3_2518 (N9372, N8466, N8463, N8480);
  not NOT1_2519 (N9375, N8497);
  not NOT1_2520 (N9381, N8766);
  not NOT1_2521 (N9382, N8778);
  not NOT1_2522 (N9383, N8793);
  not NOT1_2523 (N9384, N8796);
  and AND2_2524 (N9385, N8485, N8497);
  not NOT1_2525 (N9392, N8525);
  not NOT1_2526 (N9393, N8528);
  not NOT1_2527 (N9394, N8531);
  not NOT1_2528 (N9395, N8534);
  and AND3_2529 (N9396, N7318, N7314, N8525);
  and AND3_2530 (N9397, N8522, N8519, N8528);
  and AND3_2531 (N9398, N6131, N6127, N8531);
  and AND3_2532 (N9399, N7328, N7325, N8534);
  nor NOR2_2533 (N9400, N9024, N8539);
  nor NOR2_2534 (N9401, N9025, N8540);
  not NOT1_2535 (N9402, N8541);
  nand NAND2_2536 (N9407, N8548, N89);
  and AND2_2537 (N9408, N8541, N8548);
  not NOT1_2538 (N9412, N8811);
  not NOT1_2539 (N9413, N8566);
  not NOT1_2540 (N9414, N8569);
  not NOT1_2541 (N9415, N8572);
  not NOT1_2542 (N9416, N8575);
  nor NOR2_2543 (N9417, N9053, N8578);
  nor NOR2_2544 (N9418, N9054, N8579);
  and AND3_2545 (N9419, N7387, N6177, N8566);
  and AND3_2546 (N9420, N8555, N7384, N8569);
  and AND3_2547 (N9421, N7398, N7394, N8572);
  and AND3_2548 (N9422, N8561, N8558, N8575);
  buf BUFF1_2549 (N9423, N8326);
  nand NAND2_2550 (N9426, N9064, N8608);
  nand NAND2_2551 (N9429, N9065, N8610);
  nand NAND2_2552 (N9432, N3515, N9066);
  nand NAND2_2553 (N9435, N4796, N9072);
  nand NAND2_2554 (N9442, N3628, N9087);
  nand NAND2_2555 (N9445, N4814, N9093);
  not NOT1_2556 (N9454, N8678);
  not NOT1_2557 (N9455, N8681);
  not NOT1_2558 (N9456, N8684);
  not NOT1_2559 (N9459, N8690);
  not NOT1_2560 (N9460, N8693);
  not NOT1_2561 (N9461, N8696);
  buf BUFF1_2562 (N9462, N8358);
  not NOT1_2563 (N9465, N8702);
  not NOT1_2564 (N9466, N8705);
  not NOT1_2565 (N9467, N8708);
  not NOT1_2566 (N9468, N8724);
  buf BUFF1_2567 (N9473, N8358);
  not NOT1_2568 (N9476, N8718);
  not NOT1_2569 (N9477, N8721);
  nand NAND2_2570 (N9478, N9159, N9160);
  nand NAND2_2571 (N9485, N9179, N9180);
  nand NAND2_2572 (N9488, N9181, N9182);
  not NOT1_2573 (N9493, N8757);
  not NOT1_2574 (N9494, N8760);
  not NOT1_2575 (N9495, N8763);
  not NOT1_2576 (N9498, N8769);
  not NOT1_2577 (N9499, N8772);
  not NOT1_2578 (N9500, N8775);
  not NOT1_2579 (N9505, N8781);
  not NOT1_2580 (N9506, N8784);
  not NOT1_2581 (N9507, N8787);
  not NOT1_2582 (N9508, N8790);
  not NOT1_2583 (N9509, N8808);
  not NOT1_2584 (N9514, N8799);
  not NOT1_2585 (N9515, N8802);
  not NOT1_2586 (N9516, N8805);
  nand NAND2_2587 (N9517, N9234, N9235);
  nand NAND2_2588 (N9520, N9236, N9237);
  and AND2_2589 (N9526, N8943, N8421);
  and AND2_2590 (N9531, N8943, N8421);
  nand NAND2_2591 (N9539, N9271, N8880);
  nand NAND2_2592 (N9540, N9273, N8884);
  not NOT1_2593 (N9541, N9275);
  and AND2_2594 (N9543, N8857, N8254);
  and AND2_2595 (N9551, N8871, N8288);
  nand NAND2_2596 (N9555, N9272, N8882);
  nand NAND2_2597 (N9556, N9274, N8886);
  not NOT1_2598 (N9557, N8898);
  and AND2_2599 (N9560, N8902, N8333);
  not NOT1_2600 (N9561, N9099);
  nand NAND2_2601 (N9562, N9099, N9290);
  not NOT1_2602 (N9563, N9103);
  nand NAND2_2603 (N9564, N9103, N9292);
  not NOT1_2604 (N9565, N9107);
  nand NAND2_2605 (N9566, N9107, N9294);
  not NOT1_2606 (N9567, N9111);
  nand NAND2_2607 (N9568, N9111, N9296);
  nand NAND2_2608 (N9569, N4844, N9298);
  nand NAND2_2609 (N9570, N6207, N9300);
  not NOT1_2610 (N9571, N8920);
  not NOT1_2611 (N9575, N8927);
  and AND2_2612 (N9579, N8365, N8927);
  not NOT1_2613 (N9581, N8950);
  not NOT1_2614 (N9582, N8956);
  and AND2_2615 (N9585, N8405, N8956);
  and AND2_2616 (N9591, N8966, N8430);
  not NOT1_2617 (N9592, N9161);
  nand NAND2_2618 (N9593, N9161, N9352);
  not NOT1_2619 (N9594, N9165);
  nand NAND2_2620 (N9595, N9165, N9354);
  not NOT1_2621 (N9596, N9169);
  nand NAND2_2622 (N9597, N9169, N9356);
  not NOT1_2623 (N9598, N9173);
  nand NAND2_2624 (N9599, N9173, N9358);
  nand NAND2_2625 (N9600, N4940, N9360);
  nand NAND2_2626 (N9601, N6220, N9362);
  and AND3_2627 (N9602, N8457, N7198, N9363);
  and AND3_2628 (N9603, N7194, N8460, N9364);
  and AND3_2629 (N9604, N8463, N7209, N9365);
  and AND3_2630 (N9605, N7205, N8466, N9366);
  not NOT1_2631 (N9608, N9001);
  and AND2_2632 (N9611, N8485, N9001);
  and AND3_2633 (N9612, N8519, N7318, N9392);
  and AND3_2634 (N9613, N7314, N8522, N9393);
  and AND3_2635 (N9614, N7325, N6131, N9394);
  and AND3_2636 (N9615, N6127, N7328, N9395);
  not NOT1_2637 (N9616, N9029);
  not NOT1_2638 (N9617, N9035);
  and AND2_2639 (N9618, N8541, N9035);
  and AND3_2640 (N9621, N7384, N7387, N9413);
  and AND3_2641 (N9622, N6177, N8555, N9414);
  and AND3_2642 (N9623, N8558, N7398, N9415);
  and AND3_2643 (N9624, N7394, N8561, N9416);
  or OR5_2644 (N9626, N4563, N8352, N8353, N8354, N9285);
  or OR4_2645 (N9629, N4566, N8355, N8356, N9286);
  or OR3_2646 (N9632, N4570, N8357, N9287);
  or OR2_2647 (N9635, N5960, N9288);
  nand NAND2_2648 (N9642, N9067, N9432);
  not NOT1_2649 (N9645, N9068);
  nand NAND2_2650 (N9646, N9073, N9435);
  not NOT1_2651 (N9649, N9074);
  nand NAND2_2652 (N9650, N9257, N9256);
  nand NAND2_2653 (N9653, N9259, N9258);
  nand NAND2_2654 (N9656, N9261, N9260);
  not NOT1_2655 (N9659, N9079);
  nand NAND2_2656 (N9660, N9079, N4809);
  not NOT1_2657 (N9661, N9083);
  nand NAND2_2658 (N9662, N9083, N6202);
  nand NAND2_2659 (N9663, N9088, N9442);
  not NOT1_2660 (N9666, N9089);
  nand NAND2_2661 (N9667, N9094, N9445);
  not NOT1_2662 (N9670, N9095);
  or OR2_2663 (N9671, N8924, N8393);
  not NOT1_2664 (N9674, N9117);
  not NOT1_2665 (N9675, N8924);
  not NOT1_2666 (N9678, N9127);
  or OR4_2667 (N9679, N4597, N8388, N8389, N9315);
  or OR2_2668 (N9682, N8931, N9318);
  or OR5_2669 (N9685, N4593, N8382, N8383, N8384, N9314);
  not NOT1_2670 (N9690, N9146);
  nand NAND2_2671 (N9691, N9146, N8717);
  not NOT1_2672 (N9692, N8931);
  not NOT1_2673 (N9695, N9149);
  nand NAND2_2674 (N9698, N9401, N9400);
  nand NAND2_2675 (N9702, N9368, N9367);
  or OR2_2676 (N9707, N8996, N8517);
  not NOT1_2677 (N9710, N9183);
  not NOT1_2678 (N9711, N8996);
  not NOT1_2679 (N9714, N9193);
  not NOT1_2680 (N9715, N9203);
  nand NAND2_2681 (N9716, N9203, N6235);
  or OR2_2682 (N9717, N9005, N8518);
  not NOT1_2683 (N9720, N9206);
  not NOT1_2684 (N9721, N9220);
  nand NAND2_2685 (N9722, N9220, N7573);
  not NOT1_2686 (N9723, N9005);
  not NOT1_2687 (N9726, N9223);
  nand NAND2_2688 (N9727, N9418, N9417);
  and AND2_2689 (N9732, N9268, N8269);
  nand NAND2_2690 (N9733, N9581, N9326);
  and AND5_2691 (N9734, N89, N9408, N9332, N8394, N8421);
  and AND5_2692 (N9735, N89, N9408, N9332, N8394, N8421);
  and AND2_2693 (N9736, N9265, N8262);
  not NOT1_2694 (N9737, N9555);
  not NOT1_2695 (N9738, N9556);
  nand NAND2_2696 (N9739, N9361, N9601);
  nand NAND2_2697 (N9740, N9423, N1115);
  not NOT1_2698 (N9741, N9423);
  nand NAND2_2699 (N9742, N9299, N9570);
  and AND2_2700 (N9754, N8333, N9280);
  or OR2_2701 (N9758, N8898, N9560);
  nand NAND2_2702 (N9762, N8660, N9561);
  nand NAND2_2703 (N9763, N8663, N9563);
  nand NAND2_2704 (N9764, N8666, N9565);
  nand NAND2_2705 (N9765, N8669, N9567);
  nand NAND2_2706 (N9766, N9297, N9569);
  and AND2_2707 (N9767, N9280, N367);
  nand NAND2_2708 (N9768, N9557, N9276);
  not NOT1_2709 (N9769, N9307);
  nand NAND2_2710 (N9773, N9307, N367);
  nand NAND2_2711 (N9774, N9571, N9301);
  and AND2_2712 (N9775, N8365, N9307);
  or OR2_2713 (N9779, N8920, N9579);
  not NOT1_2714 (N9784, N9478);
  nand NAND2_2715 (N9785, N9616, N9402);
  or OR2_2716 (N9786, N8950, N9585);
  and AND4_2717 (N9790, N89, N9408, N9332, N8394);
  or OR2_2718 (N9791, N8963, N9591);
  nand NAND2_2719 (N9795, N8735, N9592);
  nand NAND2_2720 (N9796, N8738, N9594);
  nand NAND2_2721 (N9797, N8741, N9596);
  nand NAND2_2722 (N9798, N8744, N9598);
  nand NAND2_2723 (N9799, N9359, N9600);
  nor NOR2_2724 (N9800, N9602, N9369);
  nor NOR2_2725 (N9801, N9603, N9370);
  nor NOR2_2726 (N9802, N9604, N9371);
  nor NOR2_2727 (N9803, N9605, N9372);
  not NOT1_2728 (N9805, N9485);
  not NOT1_2729 (N9806, N9488);
  or OR2_2730 (N9809, N8995, N9611);
  nor NOR2_2731 (N9813, N9612, N9396);
  nor NOR2_2732 (N9814, N9613, N9397);
  nor NOR2_2733 (N9815, N9614, N9398);
  nor NOR2_2734 (N9816, N9615, N9399);
  and AND2_2735 (N9817, N9617, N9407);
  or OR2_2736 (N9820, N9029, N9618);
  not NOT1_2737 (N9825, N9517);
  not NOT1_2738 (N9826, N9520);
  nor NOR2_2739 (N9827, N9621, N9419);
  nor NOR2_2740 (N9828, N9622, N9420);
  nor NOR2_2741 (N9829, N9623, N9421);
  nor NOR2_2742 (N9830, N9624, N9422);
  not NOT1_2743 (N9835, N9426);
  nand NAND2_2744 (N9836, N9426, N4789);
  not NOT1_2745 (N9837, N9429);
  nand NAND2_2746 (N9838, N9429, N4794);
  nand NAND2_2747 (N9846, N3625, N9659);
  nand NAND2_2748 (N9847, N4810, N9661);
  not NOT1_2749 (N9862, N9462);
  nand NAND2_2750 (N9863, N7553, N9690);
  not NOT1_2751 (N9866, N9473);
  nand NAND2_2752 (N9873, N5030, N9715);
  nand NAND2_2753 (N9876, N6236, N9721);
  nand NAND2_2754 (N9890, N9795, N9593);
  nand NAND2_2755 (N9891, N9797, N9597);
  not NOT1_2756 (N9892, N9799);
  nand NAND2_2757 (N9893, N871, N9741);
  nand NAND2_2758 (N9894, N9762, N9562);
  nand NAND2_2759 (N9895, N9764, N9566);
  not NOT1_2760 (N9896, N9766);
  not NOT1_2761 (N9897, N9626);
  nand NAND2_2762 (N9898, N9626, N9249);
  not NOT1_2763 (N9899, N9629);
  nand NAND2_2764 (N9900, N9629, N9250);
  not NOT1_2765 (N9901, N9632);
  nand NAND2_2766 (N9902, N9632, N9251);
  not NOT1_2767 (N9903, N9635);
  nand NAND2_2768 (N9904, N9635, N9252);
  not NOT1_2769 (N9905, N9543);
  not NOT1_2770 (N9906, N9650);
  nand NAND2_2771 (N9907, N9650, N5769);
  not NOT1_2772 (N9908, N9653);
  nand NAND2_2773 (N9909, N9653, N5770);
  not NOT1_2774 (N9910, N9656);
  nand NAND2_2775 (N9911, N9656, N9262);
  not NOT1_2776 (N9917, N9551);
  nand NAND2_2777 (N9923, N9763, N9564);
  nand NAND2_2778 (N9924, N9765, N9568);
  or OR2_2779 (N9925, N8902, N9767);
  and AND2_2780 (N9932, N9575, N9773);
  and AND2_2781 (N9935, N9575, N9769);
  not NOT1_2782 (N9938, N9698);
  nand NAND2_2783 (N9939, N9698, N9323);
  nand NAND2_2784 (N9945, N9796, N9595);
  nand NAND2_2785 (N9946, N9798, N9599);
  not NOT1_2786 (N9947, N9702);
  nand NAND2_2787 (N9948, N9702, N6102);
  and AND2_2788 (N9949, N9608, N9375);
  not NOT1_2789 (N9953, N9727);
  nand NAND2_2790 (N9954, N9727, N9412);
  nand NAND2_2791 (N9955, N3502, N9835);
  nand NAND2_2792 (N9956, N3510, N9837);
  not NOT1_2793 (N9957, N9642);
  nand NAND2_2794 (N9958, N9642, N9645);
  not NOT1_2795 (N9959, N9646);
  nand NAND2_2796 (N9960, N9646, N9649);
  nand NAND2_2797 (N9961, N9660, N9846);
  nand NAND2_2798 (N9964, N9662, N9847);
  not NOT1_2799 (N9967, N9663);
  nand NAND2_2800 (N9968, N9663, N9666);
  not NOT1_2801 (N9969, N9667);
  nand NAND2_2802 (N9970, N9667, N9670);
  not NOT1_2803 (N9971, N9671);
  nand NAND2_2804 (N9972, N9671, N6213);
  not NOT1_2805 (N9973, N9675);
  nand NAND2_2806 (N9974, N9675, N7551);
  not NOT1_2807 (N9975, N9679);
  nand NAND2_2808 (N9976, N9679, N7552);
  not NOT1_2809 (N9977, N9682);
  not NOT1_2810 (N9978, N9685);
  nand NAND2_2811 (N9979, N9691, N9863);
  not NOT1_2812 (N9982, N9692);
  nand NAND2_2813 (N9983, N9814, N9813);
  nand NAND2_2814 (N9986, N9816, N9815);
  nand NAND2_2815 (N9989, N9801, N9800);
  nand NAND2_2816 (N9992, N9803, N9802);
  not NOT1_2817 (N9995, N9707);
  nand NAND2_2818 (N9996, N9707, N6231);
  not NOT1_2819 (N9997, N9711);
  nand NAND2_2820 (N9998, N9711, N7572);
  nand NAND2_2821 (N9999, N9716, N9873);
  not NOT1_2822 (N10002, N9717);
  nand NAND2_2823 (N10003, N9722, N9876);
  not NOT1_2824 (N10006, N9723);
  nand NAND2_2825 (N10007, N9830, N9829);
  nand NAND2_2826 (N10010, N9828, N9827);
  and AND3_2827 (N10013, N9791, N8307, N8269);
  and AND4_2828 (N10014, N9758, N9344, N8307, N8269);
  and AND5_2829 (N10015, N367, N9754, N9344, N8307, N8269);
  and AND3_2830 (N10016, N9786, N8394, N8421);
  and AND4_2831 (N10017, N9820, N9332, N8394, N8421);
  and AND3_2832 (N10018, N9786, N8394, N8421);
  and AND4_2833 (N10019, N9820, N9332, N8394, N8421);
  and AND3_2834 (N10020, N9809, N8298, N8262);
  and AND4_2835 (N10021, N9779, N9385, N8298, N8262);
  and AND5_2836 (N10022, N367, N9775, N9385, N8298, N8262);
  not NOT1_2837 (N10023, N9945);
  not NOT1_2838 (N10024, N9946);
  nand NAND2_2839 (N10025, N9740, N9893);
  not NOT1_2840 (N10026, N9923);
  not NOT1_2841 (N10028, N9924);
  nand NAND2_2842 (N10032, N8595, N9897);
  nand NAND2_2843 (N10033, N8598, N9899);
  nand NAND2_2844 (N10034, N8601, N9901);
  nand NAND2_2845 (N10035, N8604, N9903);
  nand NAND2_2846 (N10036, N4803, N9906);
  nand NAND2_2847 (N10037, N4806, N9908);
  nand NAND2_2848 (N10038, N8627, N9910);
  and AND2_2849 (N10039, N9809, N8298);
  and AND3_2850 (N10040, N9779, N9385, N8298);
  and AND4_2851 (N10041, N367, N9775, N9385, N8298);
  and AND2_2852 (N10042, N9779, N9385);
  and AND3_2853 (N10043, N367, N9775, N9385);
  nand NAND2_2854 (N10050, N8727, N9938);
  not NOT1_2855 (N10053, N9817);
  and AND2_2856 (N10054, N9817, N9029);
  and AND2_2857 (N10055, N9786, N8394);
  and AND3_2858 (N10056, N9820, N9332, N8394);
  and AND2_2859 (N10057, N9791, N8307);
  and AND3_2860 (N10058, N9758, N9344, N8307);
  and AND4_2861 (N10059, N367, N9754, N9344, N8307);
  and AND2_2862 (N10060, N9758, N9344);
  and AND3_2863 (N10061, N367, N9754, N9344);
  nand NAND2_2864 (N10062, N4997, N9947);
  nand NAND2_2865 (N10067, N8811, N9953);
  nand NAND2_2866 (N10070, N9955, N9836);
  nand NAND2_2867 (N10073, N9956, N9838);
  nand NAND2_2868 (N10076, N9068, N9957);
  nand NAND2_2869 (N10077, N9074, N9959);
  nand NAND2_2870 (N10082, N9089, N9967);
  nand NAND2_2871 (N10083, N9095, N9969);
  nand NAND2_2872 (N10084, N4871, N9971);
  nand NAND2_2873 (N10085, N6214, N9973);
  nand NAND2_2874 (N10086, N6217, N9975);
  nand NAND2_2875 (N10093, N5027, N9995);
  nand NAND2_2876 (N10094, N6232, N9997);
  or OR5_2877 (N10101, N9238, N9732, N10013, N10014, N10015);
  or OR5_2878 (N10102, N9339, N9526, N10016, N10017, N9734);
  or OR5_2879 (N10103, N9339, N9531, N10018, N10019, N9735);
  or OR5_2880 (N10104, N9242, N9736, N10020, N10021, N10022);
  and AND2_2881 (N10105, N9925, N9894);
  and AND2_2882 (N10106, N9925, N9895);
  and AND2_2883 (N10107, N9925, N9896);
  and AND2_2884 (N10108, N9925, N8253);
  nand NAND2_2885 (N10109, N10032, N9898);
  nand NAND2_2886 (N10110, N10033, N9900);
  nand NAND2_2887 (N10111, N10034, N9902);
  nand NAND2_2888 (N10112, N10035, N9904);
  nand NAND2_2889 (N10113, N10036, N9907);
  nand NAND2_2890 (N10114, N10037, N9909);
  nand NAND2_2891 (N10115, N10038, N9911);
  or OR4_2892 (N10116, N9265, N10039, N10040, N10041);
  or OR3_2893 (N10119, N9809, N10042, N10043);
  not NOT1_2894 (N10124, N9925);
  and AND2_2895 (N10130, N9768, N9925);
  not NOT1_2896 (N10131, N9932);
  not NOT1_2897 (N10132, N9935);
  and AND2_2898 (N10133, N9932, N8920);
  nand NAND2_2899 (N10134, N10050, N9939);
  not NOT1_2900 (N10135, N9983);
  nand NAND2_2901 (N10136, N9983, N9324);
  not NOT1_2902 (N10137, N9986);
  nand NAND2_2903 (N10138, N9986, N9784);
  and AND2_2904 (N10139, N9785, N10053);
  or OR4_2905 (N10140, N8943, N10055, N10056, N9790);
  or OR4_2906 (N10141, N9268, N10057, N10058, N10059);
  or OR3_2907 (N10148, N9791, N10060, N10061);
  nand NAND2_2908 (N10155, N10062, N9948);
  not NOT1_2909 (N10156, N9989);
  nand NAND2_2910 (N10157, N9989, N9805);
  not NOT1_2911 (N10158, N9992);
  nand NAND2_2912 (N10159, N9992, N9806);
  not NOT1_2913 (N10160, N9949);
  nand NAND2_2914 (N10161, N10067, N9954);
  not NOT1_2915 (N10162, N10007);
  nand NAND2_2916 (N10163, N10007, N9825);
  not NOT1_2917 (N10164, N10010);
  nand NAND2_2918 (N10165, N10010, N9826);
  nand NAND2_2919 (N10170, N10076, N9958);
  nand NAND2_2920 (N10173, N10077, N9960);
  not NOT1_2921 (N10176, N9961);
  nand NAND2_2922 (N10177, N9961, N9082);
  not NOT1_2923 (N10178, N9964);
  nand NAND2_2924 (N10179, N9964, N9086);
  nand NAND2_2925 (N10180, N10082, N9968);
  nand NAND2_2926 (N10183, N10083, N9970);
  nand NAND2_2927 (N10186, N9972, N10084);
  nand NAND2_2928 (N10189, N9974, N10085);
  nand NAND2_2929 (N10192, N9976, N10086);
  not NOT1_2930 (N10195, N9979);
  nand NAND2_2931 (N10196, N9979, N9982);
  nand NAND2_2932 (N10197, N9996, N10093);
  nand NAND2_2933 (N10200, N9998, N10094);
  not NOT1_2934 (N10203, N9999);
  nand NAND2_2935 (N10204, N9999, N10002);
  not NOT1_2936 (N10205, N10003);
  nand NAND2_2937 (N10206, N10003, N10006);
  nand NAND2_2938 (N10212, N10070, N4308);
  nand NAND2_2939 (N10213, N10073, N4313);
  and AND2_2940 (N10230, N9774, N10131);
  nand NAND2_2941 (N10231, N8730, N10135);
  nand NAND2_2942 (N10232, N9478, N10137);
  or OR2_2943 (N10233, N10139, N10054);
  nand NAND2_2944 (N10234, N7100, N10140);
  nand NAND2_2945 (N10237, N9485, N10156);
  nand NAND2_2946 (N10238, N9488, N10158);
  nand NAND2_2947 (N10239, N9517, N10162);
  nand NAND2_2948 (N10240, N9520, N10164);
  not NOT1_2949 (N10241, N10070);
  not NOT1_2950 (N10242, N10073);
  nand NAND2_2951 (N10247, N8146, N10176);
  nand NAND2_2952 (N10248, N8156, N10178);
  nand NAND2_2953 (N10259, N9692, N10195);
  nand NAND2_2954 (N10264, N9717, N10203);
  nand NAND2_2955 (N10265, N9723, N10205);
  and AND2_2956 (N10266, N10026, N10124);
  and AND2_2957 (N10267, N10028, N10124);
  and AND2_2958 (N10268, N9742, N10124);
  and AND2_2959 (N10269, N6923, N10124);
  nand NAND2_2960 (N10270, N6762, N10116);
  nand NAND2_2961 (N10271, N3061, N10241);
  nand NAND2_2962 (N10272, N3064, N10242);
  buf BUFF1_2963 (N10273, N10116);
  and AND5_2964 (N10278, N10141, N5728, N5707, N5718, N5697);
  and AND4_2965 (N10279, N10141, N5728, N5707, N5718);
  and AND3_2966 (N10280, N10141, N5728, N5718);
  and AND2_2967 (N10281, N10141, N5728);
  and AND2_2968 (N10282, N6784, N10141);
  not NOT1_2969 (N10283, N10119);
  and AND5_2970 (N10287, N10148, N5936, N5915, N5926, N5905);
  and AND4_2971 (N10288, N10148, N5936, N5915, N5926);
  and AND3_2972 (N10289, N10148, N5936, N5926);
  and AND2_2973 (N10290, N10148, N5936);
  and AND2_2974 (N10291, N6881, N10148);
  and AND2_2975 (N10292, N8898, N10124);
  nand NAND2_2976 (N10293, N10231, N10136);
  nand NAND2_2977 (N10294, N10232, N10138);
  nand NAND2_2978 (N10295, N8412, N10233);
  and AND2_2979 (N10296, N8959, N10234);
  nand NAND2_2980 (N10299, N10237, N10157);
  nand NAND2_2981 (N10300, N10238, N10159);
  or OR2_2982 (N10301, N10230, N10133);
  nand NAND2_2983 (N10306, N10239, N10163);
  nand NAND2_2984 (N10307, N10240, N10165);
  buf BUFF1_2985 (N10308, N10148);
  buf BUFF1_2986 (N10311, N10141);
  not NOT1_2987 (N10314, N10170);
  nand NAND2_2988 (N10315, N10170, N9071);
  not NOT1_2989 (N10316, N10173);
  nand NAND2_2990 (N10317, N10173, N9077);
  nand NAND2_2991 (N10318, N10247, N10177);
  nand NAND2_2992 (N10321, N10248, N10179);
  not NOT1_2993 (N10324, N10180);
  nand NAND2_2994 (N10325, N10180, N9092);
  not NOT1_2995 (N10326, N10183);
  nand NAND2_2996 (N10327, N10183, N9098);
  not NOT1_2997 (N10328, N10186);
  nand NAND2_2998 (N10329, N10186, N9674);
  not NOT1_2999 (N10330, N10189);
  nand NAND2_3000 (N10331, N10189, N9678);
  not NOT1_3001 (N10332, N10192);
  nand NAND2_3002 (N10333, N10192, N9977);
  nand NAND2_3003 (N10334, N10259, N10196);
  not NOT1_3004 (N10337, N10197);
  nand NAND2_3005 (N10338, N10197, N9710);
  not NOT1_3006 (N10339, N10200);
  nand NAND2_3007 (N10340, N10200, N9714);
  nand NAND2_3008 (N10341, N10264, N10204);
  nand NAND2_3009 (N10344, N10265, N10206);
  or OR2_3010 (N10350, N10266, N10105);
  or OR2_3011 (N10351, N10267, N10106);
  or OR2_3012 (N10352, N10268, N10107);
  or OR2_3013 (N10353, N10269, N10108);
  and AND2_3014 (N10354, N8857, N10270);
  nand NAND2_3015 (N10357, N10271, N10212);
  nand NAND2_3016 (N10360, N10272, N10213);
  or OR2_3017 (N10367, N7620, N10282);
  or OR2_3018 (N10375, N7671, N10291);
  or OR2_3019 (N10381, N10292, N10130);
  and AND4_3020 (N10388, N10114, N10134, N10293, N10294);
  and AND2_3021 (N10391, N9582, N10295);
  and AND4_3022 (N10399, N10113, N10115, N10299, N10300);
  and AND4_3023 (N10402, N10155, N10161, N10306, N10307);
  or OR5_3024 (N10406, N3229, N6888, N6889, N6890, N10287);
  or OR4_3025 (N10409, N3232, N6891, N6892, N10288);
  or OR3_3026 (N10412, N3236, N6893, N10289);
  or OR2_3027 (N10415, N3241, N10290);
  or OR5_3028 (N10419, N3137, N6791, N6792, N6793, N10278);
  or OR4_3029 (N10422, N3140, N6794, N6795, N10279);
  or OR3_3030 (N10425, N3144, N6796, N10280);
  or OR2_3031 (N10428, N3149, N10281);
  nand NAND2_3032 (N10431, N8117, N10314);
  nand NAND2_3033 (N10432, N8134, N10316);
  nand NAND2_3034 (N10437, N8169, N10324);
  nand NAND2_3035 (N10438, N8186, N10326);
  nand NAND2_3036 (N10439, N9117, N10328);
  nand NAND2_3037 (N10440, N9127, N10330);
  nand NAND2_3038 (N10441, N9682, N10332);
  nand NAND2_3039 (N10444, N9183, N10337);
  nand NAND2_3040 (N10445, N9193, N10339);
  not NOT1_3041 (N10450, N10296);
  and AND2_3042 (N10451, N10296, N4193);
  not NOT1_3043 (N10455, N10308);
  nand NAND2_3044 (N10456, N10308, N8242);
  not NOT1_3045 (N10465, N10311);
  nand NAND2_3046 (N10466, N10311, N8247);
  not NOT1_3047 (N10479, N10273);
  not NOT1_3048 (N10497, N10301);
  nand NAND2_3049 (N10509, N10431, N10315);
  nand NAND2_3050 (N10512, N10432, N10317);
  not NOT1_3051 (N10515, N10318);
  nand NAND2_3052 (N10516, N10318, N8632);
  not NOT1_3053 (N10517, N10321);
  nand NAND2_3054 (N10518, N10321, N8637);
  nand NAND2_3055 (N10519, N10437, N10325);
  nand NAND2_3056 (N10522, N10438, N10327);
  nand NAND2_3057 (N10525, N10439, N10329);
  nand NAND2_3058 (N10528, N10440, N10331);
  nand NAND2_3059 (N10531, N10441, N10333);
  not NOT1_3060 (N10534, N10334);
  nand NAND2_3061 (N10535, N10334, N9695);
  nand NAND2_3062 (N10536, N10444, N10338);
  nand NAND2_3063 (N10539, N10445, N10340);
  not NOT1_3064 (N10542, N10341);
  nand NAND2_3065 (N10543, N10341, N9720);
  not NOT1_3066 (N10544, N10344);
  nand NAND2_3067 (N10545, N10344, N9726);
  and AND2_3068 (N10546, N5631, N10450);
  not NOT1_3069 (N10547, N10391);
  and AND2_3070 (N10548, N10391, N8950);
  and AND2_3071 (N10549, N5165, N10367);
  not NOT1_3072 (N10550, N10354);
  and AND2_3073 (N10551, N10354, N3126);
  nand NAND2_3074 (N10552, N7411, N10455);
  and AND2_3075 (N10553, N10375, N9539);
  and AND2_3076 (N10554, N10375, N9540);
  and AND2_3077 (N10555, N10375, N9541);
  and AND2_3078 (N10556, N10375, N6761);
  not NOT1_3079 (N10557, N10406);
  nand NAND2_3080 (N10558, N10406, N8243);
  not NOT1_3081 (N10559, N10409);
  nand NAND2_3082 (N10560, N10409, N8244);
  not NOT1_3083 (N10561, N10412);
  nand NAND2_3084 (N10562, N10412, N8245);
  not NOT1_3085 (N10563, N10415);
  nand NAND2_3086 (N10564, N10415, N8246);
  nand NAND2_3087 (N10565, N7426, N10465);
  not NOT1_3088 (N10566, N10419);
  nand NAND2_3089 (N10567, N10419, N8248);
  not NOT1_3090 (N10568, N10422);
  nand NAND2_3091 (N10569, N10422, N8249);
  not NOT1_3092 (N10570, N10425);
  nand NAND2_3093 (N10571, N10425, N8250);
  not NOT1_3094 (N10572, N10428);
  nand NAND2_3095 (N10573, N10428, N8251);
  not NOT1_3096 (N10574, N10399);
  not NOT1_3097 (N10575, N10402);
  not NOT1_3098 (N10576, N10388);
  and AND3_3099 (N10577, N10399, N10402, N10388);
  and AND3_3100 (N10581, N10360, N9543, N10273);
  and AND3_3101 (N10582, N10357, N9905, N10273);
  not NOT1_3102 (N10583, N10367);
  and AND2_3103 (N10587, N10367, N5735);
  and AND2_3104 (N10588, N10367, N3135);
  not NOT1_3105 (N10589, N10375);
  and AND5_3106 (N10594, N10381, N7180, N7159, N7170, N7149);
  and AND4_3107 (N10595, N10381, N7180, N7159, N7170);
  and AND3_3108 (N10596, N10381, N7180, N7170);
  and AND2_3109 (N10597, N10381, N7180);
  and AND2_3110 (N10598, N8444, N10381);
  buf BUFF1_3111 (N10602, N10381);
  nand NAND2_3112 (N10609, N7479, N10515);
  nand NAND2_3113 (N10610, N7491, N10517);
  nand NAND2_3114 (N10621, N9149, N10534);
  nand NAND2_3115 (N10626, N9206, N10542);
  nand NAND2_3116 (N10627, N9223, N10544);
  or OR2_3117 (N10628, N10546, N10451);
  and AND2_3118 (N10629, N9733, N10547);
  and AND2_3119 (N10631, N5166, N10550);
  nand NAND2_3120 (N10632, N10552, N10456);
  nand NAND2_3121 (N10637, N7414, N10557);
  nand NAND2_3122 (N10638, N7417, N10559);
  nand NAND2_3123 (N10639, N7420, N10561);
  nand NAND2_3124 (N10640, N7423, N10563);
  nand NAND2_3125 (N10641, N10565, N10466);
  nand NAND2_3126 (N10642, N7429, N10566);
  nand NAND2_3127 (N10643, N7432, N10568);
  nand NAND2_3128 (N10644, N7435, N10570);
  nand NAND2_3129 (N10645, N7438, N10572);
  and AND3_3130 (N10647, N886, N887, N10577);
  and AND3_3131 (N10648, N10360, N8857, N10479);
  and AND3_3132 (N10649, N10357, N7609, N10479);
  or OR2_3133 (N10652, N8966, N10598);
  or OR5_3134 (N10659, N4675, N8451, N8452, N8453, N10594);
  or OR4_3135 (N10662, N4678, N8454, N8455, N10595);
  or OR3_3136 (N10665, N4682, N8456, N10596);
  or OR2_3137 (N10668, N4687, N10597);
  not NOT1_3138 (N10671, N10509);
  nand NAND2_3139 (N10672, N10509, N8615);
  not NOT1_3140 (N10673, N10512);
  nand NAND2_3141 (N10674, N10512, N8624);
  nand NAND2_3142 (N10675, N10609, N10516);
  nand NAND2_3143 (N10678, N10610, N10518);
  not NOT1_3144 (N10681, N10519);
  nand NAND2_3145 (N10682, N10519, N8644);
  not NOT1_3146 (N10683, N10522);
  nand NAND2_3147 (N10684, N10522, N8653);
  not NOT1_3148 (N10685, N10525);
  nand NAND2_3149 (N10686, N10525, N9454);
  not NOT1_3150 (N10687, N10528);
  nand NAND2_3151 (N10688, N10528, N9459);
  not NOT1_3152 (N10689, N10531);
  nand NAND2_3153 (N10690, N10531, N9978);
  nand NAND2_3154 (N10691, N10621, N10535);
  not NOT1_3155 (N10694, N10536);
  nand NAND2_3156 (N10695, N10536, N9493);
  not NOT1_3157 (N10696, N10539);
  nand NAND2_3158 (N10697, N10539, N9498);
  nand NAND2_3159 (N10698, N10626, N10543);
  nand NAND2_3160 (N10701, N10627, N10545);
  or OR2_3161 (N10704, N10629, N10548);
  and AND2_3162 (N10705, N3159, N10583);
  or OR2_3163 (N10706, N10631, N10551);
  and AND2_3164 (N10707, N9737, N10589);
  and AND2_3165 (N10708, N9738, N10589);
  and AND2_3166 (N10709, N9243, N10589);
  and AND2_3167 (N10710, N5892, N10589);
  nand NAND2_3168 (N10711, N10637, N10558);
  nand NAND2_3169 (N10712, N10638, N10560);
  nand NAND2_3170 (N10713, N10639, N10562);
  nand NAND2_3171 (N10714, N10640, N10564);
  nand NAND2_3172 (N10715, N10642, N10567);
  nand NAND2_3173 (N10716, N10643, N10569);
  nand NAND2_3174 (N10717, N10644, N10571);
  nand NAND2_3175 (N10718, N10645, N10573);
  not NOT1_3176 (N10719, N10602);
  nand NAND2_3177 (N10720, N10602, N9244);
  not NOT1_3178 (N10729, N10647);
  and AND2_3179 (N10730, N5178, N10583);
  and AND2_3180 (N10731, N2533, N10583);
  nand NAND2_3181 (N10737, N7447, N10671);
  nand NAND2_3182 (N10738, N7465, N10673);
  or OR4_3183 (N10739, N10648, N10649, N10581, N10582);
  nand NAND2_3184 (N10746, N7503, N10681);
  nand NAND2_3185 (N10747, N7521, N10683);
  nand NAND2_3186 (N10748, N8678, N10685);
  nand NAND2_3187 (N10749, N8690, N10687);
  nand NAND2_3188 (N10750, N9685, N10689);
  nand NAND2_3189 (N10753, N8757, N10694);
  nand NAND2_3190 (N10754, N8769, N10696);
  or OR2_3191 (N10759, N10705, N10549);
  or OR2_3192 (N10760, N10707, N10553);
  or OR2_3193 (N10761, N10708, N10554);
  or OR2_3194 (N10762, N10709, N10555);
  or OR2_3195 (N10763, N10710, N10556);
  nand NAND2_3196 (N10764, N8580, N10719);
  and AND2_3197 (N10765, N10652, N9890);
  and AND2_3198 (N10766, N10652, N9891);
  and AND2_3199 (N10767, N10652, N9892);
  and AND2_3200 (N10768, N10652, N8252);
  not NOT1_3201 (N10769, N10659);
  nand NAND2_3202 (N10770, N10659, N9245);
  not NOT1_3203 (N10771, N10662);
  nand NAND2_3204 (N10772, N10662, N9246);
  not NOT1_3205 (N10773, N10665);
  nand NAND2_3206 (N10774, N10665, N9247);
  not NOT1_3207 (N10775, N10668);
  nand NAND2_3208 (N10776, N10668, N9248);
  or OR2_3209 (N10778, N10730, N10587);
  or OR2_3210 (N10781, N10731, N10588);
  not NOT1_3211 (N10784, N10652);
  nand NAND2_3212 (N10789, N10737, N10672);
  nand NAND2_3213 (N10792, N10738, N10674);
  not NOT1_3214 (N10796, N10675);
  nand NAND2_3215 (N10797, N10675, N8633);
  not NOT1_3216 (N10798, N10678);
  nand NAND2_3217 (N10799, N10678, N8638);
  nand NAND2_3218 (N10800, N10746, N10682);
  nand NAND2_3219 (N10803, N10747, N10684);
  nand NAND2_3220 (N10806, N10748, N10686);
  nand NAND2_3221 (N10809, N10749, N10688);
  nand NAND2_3222 (N10812, N10750, N10690);
  not NOT1_3223 (N10815, N10691);
  nand NAND2_3224 (N10816, N10691, N9866);
  nand NAND2_3225 (N10817, N10753, N10695);
  nand NAND2_3226 (N10820, N10754, N10697);
  not NOT1_3227 (N10823, N10698);
  nand NAND2_3228 (N10824, N10698, N9505);
  not NOT1_3229 (N10825, N10701);
  nand NAND2_3230 (N10826, N10701, N9514);
  nand NAND2_3231 (N10827, N10764, N10720);
  nand NAND2_3232 (N10832, N8583, N10769);
  nand NAND2_3233 (N10833, N8586, N10771);
  nand NAND2_3234 (N10834, N8589, N10773);
  nand NAND2_3235 (N10835, N8592, N10775);
  not NOT1_3236 (N10836, N10739);
  buf BUFF1_3237 (N10837, N10778);
  buf BUFF1_3238 (N10838, N10778);
  buf BUFF1_3239 (N10839, N10781);
  buf BUFF1_3240 (N10840, N10781);
  nand NAND2_3241 (N10845, N7482, N10796);
  nand NAND2_3242 (N10846, N7494, N10798);
  nand NAND2_3243 (N10857, N9473, N10815);
  nand NAND2_3244 (N10862, N8781, N10823);
  nand NAND2_3245 (N10863, N8799, N10825);
  and AND2_3246 (N10864, N10023, N10784);
  and AND2_3247 (N10865, N10024, N10784);
  and AND2_3248 (N10866, N9739, N10784);
  and AND2_3249 (N10867, N7136, N10784);
  nand NAND2_3250 (N10868, N10832, N10770);
  nand NAND2_3251 (N10869, N10833, N10772);
  nand NAND2_3252 (N10870, N10834, N10774);
  nand NAND2_3253 (N10871, N10835, N10776);
  not NOT1_3254 (N10872, N10789);
  nand NAND2_3255 (N10873, N10789, N8616);
  not NOT1_3256 (N10874, N10792);
  nand NAND2_3257 (N10875, N10792, N8625);
  nand NAND2_3258 (N10876, N10845, N10797);
  nand NAND2_3259 (N10879, N10846, N10799);
  not NOT1_3260 (N10882, N10800);
  nand NAND2_3261 (N10883, N10800, N8645);
  not NOT1_3262 (N10884, N10803);
  nand NAND2_3263 (N10885, N10803, N8654);
  not NOT1_3264 (N10886, N10806);
  nand NAND2_3265 (N10887, N10806, N9455);
  not NOT1_3266 (N10888, N10809);
  nand NAND2_3267 (N10889, N10809, N9460);
  not NOT1_3268 (N10890, N10812);
  nand NAND2_3269 (N10891, N10812, N9862);
  nand NAND2_3270 (N10892, N10857, N10816);
  not NOT1_3271 (N10895, N10817);
  nand NAND2_3272 (N10896, N10817, N9494);
  not NOT1_3273 (N10897, N10820);
  nand NAND2_3274 (N10898, N10820, N9499);
  nand NAND2_3275 (N10899, N10862, N10824);
  nand NAND2_3276 (N10902, N10863, N10826);
  or OR2_3277 (N10905, N10864, N10765);
  or OR2_3278 (N10906, N10865, N10766);
  or OR2_3279 (N10907, N10866, N10767);
  or OR2_3280 (N10908, N10867, N10768);
  nand NAND2_3281 (N10909, N7450, N10872);
  nand NAND2_3282 (N10910, N7468, N10874);
  nand NAND2_3283 (N10915, N7506, N10882);
  nand NAND2_3284 (N10916, N7524, N10884);
  nand NAND2_3285 (N10917, N8681, N10886);
  nand NAND2_3286 (N10918, N8693, N10888);
  nand NAND2_3287 (N10919, N9462, N10890);
  nand NAND2_3288 (N10922, N8760, N10895);
  nand NAND2_3289 (N10923, N8772, N10897);
  nand NAND2_3290 (N10928, N10909, N10873);
  nand NAND2_3291 (N10931, N10910, N10875);
  not NOT1_3292 (N10934, N10876);
  nand NAND2_3293 (N10935, N10876, N8634);
  not NOT1_3294 (N10936, N10879);
  nand NAND2_3295 (N10937, N10879, N8639);
  nand NAND2_3296 (N10938, N10915, N10883);
  nand NAND2_3297 (N10941, N10916, N10885);
  nand NAND2_3298 (N10944, N10917, N10887);
  nand NAND2_3299 (N10947, N10918, N10889);
  nand NAND2_3300 (N10950, N10919, N10891);
  not NOT1_3301 (N10953, N10892);
  nand NAND2_3302 (N10954, N10892, N9476);
  nand NAND2_3303 (N10955, N10922, N10896);
  nand NAND2_3304 (N10958, N10923, N10898);
  not NOT1_3305 (N10961, N10899);
  nand NAND2_3306 (N10962, N10899, N9506);
  not NOT1_3307 (N10963, N10902);
  nand NAND2_3308 (N10964, N10902, N9515);
  nand NAND2_3309 (N10969, N7485, N10934);
  nand NAND2_3310 (N10970, N7497, N10936);
  nand NAND2_3311 (N10981, N8718, N10953);
  nand NAND2_3312 (N10986, N8784, N10961);
  nand NAND2_3313 (N10987, N8802, N10963);
  not NOT1_3314 (N10988, N10928);
  nand NAND2_3315 (N10989, N10928, N8617);
  not NOT1_3316 (N10990, N10931);
  nand NAND2_3317 (N10991, N10931, N8626);
  nand NAND2_3318 (N10992, N10969, N10935);
  nand NAND2_3319 (N10995, N10970, N10937);
  not NOT1_3320 (N10998, N10938);
  nand NAND2_3321 (N10999, N10938, N8646);
  not NOT1_3322 (N11000, N10941);
  nand NAND2_3323 (N11001, N10941, N8655);
  not NOT1_3324 (N11002, N10944);
  nand NAND2_3325 (N11003, N10944, N9456);
  not NOT1_3326 (N11004, N10947);
  nand NAND2_3327 (N11005, N10947, N9461);
  not NOT1_3328 (N11006, N10950);
  nand NAND2_3329 (N11007, N10950, N9465);
  nand NAND2_3330 (N11008, N10981, N10954);
  not NOT1_3331 (N11011, N10955);
  nand NAND2_3332 (N11012, N10955, N9495);
  not NOT1_3333 (N11013, N10958);
  nand NAND2_3334 (N11014, N10958, N9500);
  nand NAND2_3335 (N11015, N10986, N10962);
  nand NAND2_3336 (N11018, N10987, N10964);
  nand NAND2_3337 (N11023, N7453, N10988);
  nand NAND2_3338 (N11024, N7471, N10990);
  nand NAND2_3339 (N11027, N7509, N10998);
  nand NAND2_3340 (N11028, N7527, N11000);
  nand NAND2_3341 (N11029, N8684, N11002);
  nand NAND2_3342 (N11030, N8696, N11004);
  nand NAND2_3343 (N11031, N8702, N11006);
  nand NAND2_3344 (N11034, N8763, N11011);
  nand NAND2_3345 (N11035, N8775, N11013);
  not NOT1_3346 (N11040, N10992);
  nand NAND2_3347 (N11041, N10992, N8294);
  not NOT1_3348 (N11042, N10995);
  nand NAND2_3349 (N11043, N10995, N8295);
  nand NAND2_3350 (N11044, N11023, N10989);
  nand NAND2_3351 (N11047, N11024, N10991);
  nand NAND2_3352 (N11050, N11027, N10999);
  nand NAND2_3353 (N11053, N11028, N11001);
  nand NAND2_3354 (N11056, N11029, N11003);
  nand NAND2_3355 (N11059, N11030, N11005);
  nand NAND2_3356 (N11062, N11031, N11007);
  not NOT1_3357 (N11065, N11008);
  nand NAND2_3358 (N11066, N11008, N9477);
  nand NAND2_3359 (N11067, N11034, N11012);
  nand NAND2_3360 (N11070, N11035, N11014);
  not NOT1_3361 (N11073, N11015);
  nand NAND2_3362 (N11074, N11015, N9507);
  not NOT1_3363 (N11075, N11018);
  nand NAND2_3364 (N11076, N11018, N9516);
  nand NAND2_3365 (N11077, N7488, N11040);
  nand NAND2_3366 (N11078, N7500, N11042);
  nand NAND2_3367 (N11095, N8721, N11065);
  nand NAND2_3368 (N11098, N8787, N11073);
  nand NAND2_3369 (N11099, N8805, N11075);
  nand NAND2_3370 (N11100, N11077, N11041);
  nand NAND2_3371 (N11103, N11078, N11043);
  not NOT1_3372 (N11106, N11056);
  nand NAND2_3373 (N11107, N11056, N9319);
  not NOT1_3374 (N11108, N11059);
  nand NAND2_3375 (N11109, N11059, N9320);
  not NOT1_3376 (N11110, N11067);
  nand NAND2_3377 (N11111, N11067, N9381);
  not NOT1_3378 (N11112, N11070);
  nand NAND2_3379 (N11113, N11070, N9382);
  not NOT1_3380 (N11114, N11044);
  nand NAND2_3381 (N11115, N11044, N8618);
  not NOT1_3382 (N11116, N11047);
  nand NAND2_3383 (N11117, N11047, N8619);
  not NOT1_3384 (N11118, N11050);
  nand NAND2_3385 (N11119, N11050, N8647);
  not NOT1_3386 (N11120, N11053);
  nand NAND2_3387 (N11121, N11053, N8648);
  not NOT1_3388 (N11122, N11062);
  nand NAND2_3389 (N11123, N11062, N9466);
  nand NAND2_3390 (N11124, N11095, N11066);
  nand NAND2_3391 (N11127, N11098, N11074);
  nand NAND2_3392 (N11130, N11099, N11076);
  nand NAND2_3393 (N11137, N8687, N11106);
  nand NAND2_3394 (N11138, N8699, N11108);
  nand NAND2_3395 (N11139, N8766, N11110);
  nand NAND2_3396 (N11140, N8778, N11112);
  nand NAND2_3397 (N11141, N7456, N11114);
  nand NAND2_3398 (N11142, N7474, N11116);
  nand NAND2_3399 (N11143, N7512, N11118);
  nand NAND2_3400 (N11144, N7530, N11120);
  nand NAND2_3401 (N11145, N8705, N11122);
  and AND3_3402 (N11152, N11103, N8871, N10283);
  and AND3_3403 (N11153, N11100, N7655, N10283);
  and AND3_3404 (N11154, N11103, N9551, N10119);
  and AND3_3405 (N11155, N11100, N9917, N10119);
  nand NAND2_3406 (N11156, N11137, N11107);
  nand NAND2_3407 (N11159, N11138, N11109);
  nand NAND2_3408 (N11162, N11139, N11111);
  nand NAND2_3409 (N11165, N11140, N11113);
  nand NAND2_3410 (N11168, N11141, N11115);
  nand NAND2_3411 (N11171, N11142, N11117);
  nand NAND2_3412 (N11174, N11143, N11119);
  nand NAND2_3413 (N11177, N11144, N11121);
  nand NAND2_3414 (N11180, N11145, N11123);
  not NOT1_3415 (N11183, N11124);
  nand NAND2_3416 (N11184, N11124, N9468);
  not NOT1_3417 (N11185, N11127);
  nand NAND2_3418 (N11186, N11127, N9508);
  not NOT1_3419 (N11187, N11130);
  nand NAND2_3420 (N11188, N11130, N9509);
  or OR4_3421 (N11205, N11152, N11153, N11154, N11155);
  nand NAND2_3422 (N11210, N8724, N11183);
  nand NAND2_3423 (N11211, N8790, N11185);
  nand NAND2_3424 (N11212, N8808, N11187);
  not NOT1_3425 (N11213, N11168);
  nand NAND2_3426 (N11214, N11168, N8260);
  not NOT1_3427 (N11215, N11171);
  nand NAND2_3428 (N11216, N11171, N8261);
  not NOT1_3429 (N11217, N11174);
  nand NAND2_3430 (N11218, N11174, N8296);
  not NOT1_3431 (N11219, N11177);
  nand NAND2_3432 (N11220, N11177, N8297);
  and AND3_3433 (N11222, N11159, N9575, N1218);
  and AND3_3434 (N11223, N11156, N8927, N1218);
  and AND3_3435 (N11224, N11159, N9935, N750);
  and AND3_3436 (N11225, N11156, N10132, N750);
  and AND3_3437 (N11226, N11165, N9608, N10497);
  and AND3_3438 (N11227, N11162, N9001, N10497);
  and AND3_3439 (N11228, N11165, N9949, N10301);
  and AND3_3440 (N11229, N11162, N10160, N10301);
  not NOT1_3441 (N11231, N11180);
  nand NAND2_3442 (N11232, N11180, N9467);
  nand NAND2_3443 (N11233, N11210, N11184);
  nand NAND2_3444 (N11236, N11211, N11186);
  nand NAND2_3445 (N11239, N11212, N11188);
  nand NAND2_3446 (N11242, N7459, N11213);
  nand NAND2_3447 (N11243, N7462, N11215);
  nand NAND2_3448 (N11244, N7515, N11217);
  nand NAND2_3449 (N11245, N7518, N11219);
  not NOT1_3450 (N11246, N11205);
  nand NAND2_3451 (N11250, N8708, N11231);
  or OR4_3452 (N11252, N11222, N11223, N11224, N11225);
  or OR4_3453 (N11257, N11226, N11227, N11228, N11229);
  nand NAND2_3454 (N11260, N11242, N11214);
  nand NAND2_3455 (N11261, N11243, N11216);
  nand NAND2_3456 (N11262, N11244, N11218);
  nand NAND2_3457 (N11263, N11245, N11220);
  not NOT1_3458 (N11264, N11233);
  nand NAND2_3459 (N11265, N11233, N9322);
  not NOT1_3460 (N11267, N11236);
  nand NAND2_3461 (N11268, N11236, N9383);
  not NOT1_3462 (N11269, N11239);
  nand NAND2_3463 (N11270, N11239, N9384);
  nand NAND2_3464 (N11272, N11250, N11232);
  not NOT1_3465 (N11277, N11261);
  and AND2_3466 (N11278, N10273, N11260);
  not NOT1_3467 (N11279, N11263);
  and AND2_3468 (N11280, N10119, N11262);
  nand NAND2_3469 (N11282, N8714, N11264);
  not NOT1_3470 (N11283, N11252);
  nand NAND2_3471 (N11284, N8793, N11267);
  nand NAND2_3472 (N11285, N8796, N11269);
  not NOT1_3473 (N11286, N11257);
  and AND2_3474 (N11288, N11277, N10479);
  and AND2_3475 (N11289, N11279, N10283);
  not NOT1_3476 (N11290, N11272);
  nand NAND2_3477 (N11291, N11272, N9321);
  nand NAND2_3478 (N11292, N11282, N11265);
  nand NAND2_3479 (N11293, N11284, N11268);
  nand NAND2_3480 (N11294, N11285, N11270);
  nand NAND2_3481 (N11295, N8711, N11290);
  not NOT1_3482 (N11296, N11292);
  not NOT1_3483 (N11297, N11294);
  and AND2_3484 (N11298, N10301, N11293);
  or OR2_3485 (N11299, N11288, N11278);
  or OR2_3486 (N11302, N11289, N11280);
  nand NAND2_3487 (N11307, N11295, N11291);
  and AND2_3488 (N11308, N11296, N1218);
  and AND2_3489 (N11309, N11297, N10497);
  nand NAND2_3490 (N11312, N11302, N11246);
  nand NAND2_3491 (N11313, N11299, N10836);
  not NOT1_3492 (N11314, N11299);
  not NOT1_3493 (N11315, N11302);
  and AND2_3494 (N11316, N750, N11307);
  or OR2_3495 (N11317, N11309, N11298);
  nand NAND2_3496 (N11320, N11205, N11315);
  nand NAND2_3497 (N11321, N10739, N11314);
  or OR2_3498 (N11323, N11308, N11316);
  nand NAND2_3499 (N11327, N11312, N11320);
  nand NAND2_3500 (N11328, N11313, N11321);
  nand NAND2_3501 (N11329, N11317, N11286);
  not NOT1_3502 (N11331, N11317);
  not NOT1_3503 (N11333, N11327);
  not NOT1_3504 (N11334, N11328);
  nand NAND2_3505 (N11335, N11257, N11331);
  nand NAND2_3506 (N11336, N11323, N11283);
  not NOT1_3507 (N11337, N11323);
  nand NAND2_3508 (N11338, N11329, N11335);
  nand NAND2_3509 (N11339, N11252, N11337);
  not NOT1_3510 (N11340, N11338);
  nand NAND2_3511 (N11341, N11336, N11339);
  not NOT1_3512 (N11342, N11341);
  buf BUFF1_3513 (N241_O, N241_I);

endmodule
