// AES sbox - Converted from Usuba outputs
// deyuan, 05/19/2025

module aes_sbox_usuba (
    input  wire [7:0] A,
    output wire [7:0] S
);

wire y14__ = A[4] ^ A[2];
wire y13__ = A[7] ^ A[1];
wire y9__  = A[7] ^ A[4];
wire y8__  = A[7] ^ A[2];
wire t0__  = A[6] ^ A[5];
wire y12__ = y13__ ^ y14__;
wire y1__  = t0__ ^ A[0];
wire t1__  = A[3] ^ y12__;
wire y4__  = y1__ ^ A[4];
wire y2__  = y1__ ^ A[7];
wire y5__  = y1__ ^ A[1];
wire y15__ = t1__ ^ A[2];
wire y20__ = t1__ ^ A[6];
wire t5__  = y4__ & A[0];
wire y3__  = y5__ ^ y8__;
wire t8__  = y5__ & y1__;
wire y6__  = y15__ ^ A[0];
wire y10__ = y15__ ^ t0__;
wire t2__  = y12__ & y15__;
wire y11__ = y20__ ^ y9__;
wire t3__  = y3__ & y6__;
wire y19__ = y10__ ^ y8__;
wire t15__ = y8__ & y10__;
wire t6__  = t5__ ^ t2__;
wire y7__  = A[0] ^ y11__;
wire y17__ = y10__ ^ y11__;
wire y16__ = t0__ ^ y11__;
wire t12__ = y9__ & y11__;
wire t4__  = t3__ ^ t2__;
wire t10__ = y2__ & y7__;
wire t13__ = y14__ & y17__;
wire y21__ = y13__ ^ y16__;
wire y18__ = A[7] ^ y16__;
wire t7__  = y13__ & y16__;
wire t16__ = t15__ ^ t12__;
wire t17__ = t4__ ^ y20__;
wire t14__ = t13__ ^ t12__;
wire t9__  = t8__ ^ t7__;
wire t11__ = t10__ ^ t7__;
wire t18__ = t6__ ^ t16__;
wire t21__ = t17__ ^ t14__;
wire t19__ = t9__ ^ t14__;
wire t20__ = t11__ ^ t16__;
wire t22__ = t18__ ^ y19__;
wire t23__ = t19__ ^ y21__;
wire t24__ = t20__ ^ y18__;
wire t25__ = t21__ ^ t22__;
wire t26__ = t21__ & t23__;
wire t30__ = t23__ ^ t24__;
wire t27__ = t24__ ^ t26__;
wire t31__ = t22__ ^ t26__;
wire t28__ = t25__ & t27__;
wire t32__ = t31__ & t30__;
wire t29__ = t28__ ^ t22__;
wire t33__ = t32__ ^ t24__;
wire z5__  = t29__ & y7__;
wire z14__ = t29__ & y2__;
wire t34__ = t23__ ^ t33__;
wire t35__ = t27__ ^ t33__;
wire t42__ = t29__ ^ t33__;
wire z2__  = t33__ & A[0];
wire z11__ = t33__ & y4__;
wire t36__ = t24__ & t35__;
wire z6__  = t42__ & y11__;
wire z15__ = t42__ & y9__;
wire t37__ = t36__ ^ t34__;
wire t38__ = t27__ ^ t36__;
wire t44__ = t33__ ^ t37__;
wire z1__  = t37__ & y6__;
wire z10__ = t37__ & y3__;
wire t39__ = t29__ & t38__;
wire z0__  = t44__ & y15__;
wire z9__  = t44__ & y12__;
wire t40__ = t25__ ^ t39__;
wire tc4__  = z0__ ^ z2__;
wire tc5__  = z1__ ^ z0__;
wire t41__  = t40__ ^ t37__;
wire t43__  = t29__ ^ t40__;
wire z4__   = t40__ & y1__;
wire z13__  = t40__ & y5__;
wire t45__  = t42__ ^ t41__;
wire z8__   = t41__ & y10__;
wire z17__  = t41__ & y8__;
wire z3__   = t43__ & y16__;
wire z12__  = t43__ & y13__;
wire z7__   = t45__ & y17__;
wire z16__  = t45__ & y14__;
wire tc6__  = z3__ ^ z4__;
wire tc12__ = z3__ ^ z5__;
wire tc7__  = z12__ ^ tc4__;
wire tc1__  = z15__ ^ z16__;
wire tc8__  = z7__ ^ tc6__;
wire tc11__ = tc6__ ^ tc5__;
wire tc14__ = tc4__ ^ tc12__;
wire tc9__  = z8__ ^ tc7__;
wire tc2__  = z10__ ^ tc1__;
wire tc13__ = z13__ ^ tc1__;
wire tc16__ = z6__ ^ tc8__;
wire tc10__ = tc8__ ^ tc9__;
wire tc3__  = z9__ ^ tc2__;
wire tc21__ = tc2__ ^ z11__;
wire tc18__ = tc13__ ^ tc14__;
wire tc20__ = z15__ ^ tc16__;
wire tc17__ = z14__ ^ tc10__;
wire S3__   = tc3__ ^ tc11__;
wire S0__   = tc3__ ^ tc16__;
wire _tmp1_ = z12__ ^ tc18__;
wire _tmp2_ = tc10__ ^ tc18__;
wire tc26__ = tc17__ ^ tc20__;
wire S5__   = tc21__ ^ tc17__;
wire S4__   = tc14__ ^ S3__;
wire _tmp3_ = S3__ ^ tc16__;
wire S7__   = ~_tmp1_;
wire S6__   = ~_tmp2_;
wire _tmp4_ = tc26__ ^ z17__;
wire S1__   = ~_tmp3_;
wire S2__   = ~_tmp4_;

assign S[7] = S0__;
assign S[6] = S1__;
assign S[5] = S2__;
assign S[4] = S3__;
assign S[3] = S4__;
assign S[2] = S5__;
assign S[1] = S6__;
assign S[0] = S7__;

endmodule

