// AES inverse S-box
// hosein, 03/28/2025

module aes_inverse_sbox(
    input  [7:0] pi0,
    output [7:0] po0
);

assign po0 =
    (pi0 == 8'h00) ? 8'h52 :
    (pi0 == 8'h01) ? 8'h09 :
    (pi0 == 8'h02) ? 8'h6A :
    (pi0 == 8'h03) ? 8'hD5 :
    (pi0 == 8'h04) ? 8'h30 :
    (pi0 == 8'h05) ? 8'h36 :
    (pi0 == 8'h06) ? 8'hA5 :
    (pi0 == 8'h07) ? 8'h38 :
    (pi0 == 8'h08) ? 8'hBF :
    (pi0 == 8'h09) ? 8'h40 :
    (pi0 == 8'h0A) ? 8'hA3 :
    (pi0 == 8'h0B) ? 8'h9E :
    (pi0 == 8'h0C) ? 8'h81 :
    (pi0 == 8'h0D) ? 8'hF3 :
    (pi0 == 8'h0E) ? 8'hD7 :
    (pi0 == 8'h0F) ? 8'hFB :
    (pi0 == 8'h10) ? 8'h7C :
    (pi0 == 8'h11) ? 8'hE3 :
    (pi0 == 8'h12) ? 8'h39 :
    (pi0 == 8'h13) ? 8'h82 :
    (pi0 == 8'h14) ? 8'h9B :
    (pi0 == 8'h15) ? 8'h2F :
    (pi0 == 8'h16) ? 8'hFF :
    (pi0 == 8'h17) ? 8'h87 :
    (pi0 == 8'h18) ? 8'h34 :
    (pi0 == 8'h19) ? 8'h8E :
    (pi0 == 8'h1A) ? 8'h43 :
    (pi0 == 8'h1B) ? 8'h44 :
    (pi0 == 8'h1C) ? 8'hC4 :
    (pi0 == 8'h1D) ? 8'hDE :
    (pi0 == 8'h1E) ? 8'hE9 :
    (pi0 == 8'h1F) ? 8'hCB :
    (pi0 == 8'h20) ? 8'h54 :
    (pi0 == 8'h21) ? 8'h7B :
    (pi0 == 8'h22) ? 8'h94 :
    (pi0 == 8'h23) ? 8'h32 :
    (pi0 == 8'h24) ? 8'hA6 :
    (pi0 == 8'h25) ? 8'hC2 :
    (pi0 == 8'h26) ? 8'h23 :
    (pi0 == 8'h27) ? 8'h3D :
    (pi0 == 8'h28) ? 8'hEE :
    (pi0 == 8'h29) ? 8'h4C :
    (pi0 == 8'h2A) ? 8'h95 :
    (pi0 == 8'h2B) ? 8'h0B :
    (pi0 == 8'h2C) ? 8'h42 :
    (pi0 == 8'h2D) ? 8'hFA :
    (pi0 == 8'h2E) ? 8'hC3 :
    (pi0 == 8'h2F) ? 8'h4E :
    (pi0 == 8'h30) ? 8'h08 :
    (pi0 == 8'h31) ? 8'h2E :
    (pi0 == 8'h32) ? 8'hA1 :
    (pi0 == 8'h33) ? 8'h66 :
    (pi0 == 8'h34) ? 8'h28 :
    (pi0 == 8'h35) ? 8'hD9 :
    (pi0 == 8'h36) ? 8'h24 :
    (pi0 == 8'h37) ? 8'hB2 :
    (pi0 == 8'h38) ? 8'h76 :
    (pi0 == 8'h39) ? 8'h5B :
    (pi0 == 8'h3A) ? 8'hA2 :
    (pi0 == 8'h3B) ? 8'h49 :
    (pi0 == 8'h3C) ? 8'h6D :
    (pi0 == 8'h3D) ? 8'h8B :
    (pi0 == 8'h3E) ? 8'hD1 :
    (pi0 == 8'h3F) ? 8'h25 :
    (pi0 == 8'h40) ? 8'h72 :
    (pi0 == 8'h41) ? 8'hF8 :
    (pi0 == 8'h42) ? 8'hF6 :
    (pi0 == 8'h43) ? 8'h64 :
    (pi0 == 8'h44) ? 8'h86 :
    (pi0 == 8'h45) ? 8'h68 :
    (pi0 == 8'h46) ? 8'h98 :
    (pi0 == 8'h47) ? 8'h16 :
    (pi0 == 8'h48) ? 8'hD4 :
    (pi0 == 8'h49) ? 8'hA4 :
    (pi0 == 8'h4A) ? 8'h5C :
    (pi0 == 8'h4B) ? 8'hCC :
    (pi0 == 8'h4C) ? 8'h5D :
    (pi0 == 8'h4D) ? 8'h65 :
    (pi0 == 8'h4E) ? 8'hB6 :
    (pi0 == 8'h4F) ? 8'h92 :
    (pi0 == 8'h50) ? 8'h6C :
    (pi0 == 8'h51) ? 8'h70 :
    (pi0 == 8'h52) ? 8'h48 :
    (pi0 == 8'h53) ? 8'h50 :
    (pi0 == 8'h54) ? 8'hFD :
    (pi0 == 8'h55) ? 8'hED :
    (pi0 == 8'h56) ? 8'hB9 :
    (pi0 == 8'h57) ? 8'hDA :
    (pi0 == 8'h58) ? 8'h5E :
    (pi0 == 8'h59) ? 8'h15 :
    (pi0 == 8'h5A) ? 8'h46 :
    (pi0 == 8'h5B) ? 8'h57 :
    (pi0 == 8'h5C) ? 8'hA7 :
    (pi0 == 8'h5D) ? 8'h8D :
    (pi0 == 8'h5E) ? 8'h9D :
    (pi0 == 8'h5F) ? 8'h84 :
    (pi0 == 8'h60) ? 8'h90 :
    (pi0 == 8'h61) ? 8'hD8 :
    (pi0 == 8'h62) ? 8'hAB :
    (pi0 == 8'h63) ? 8'h00 :
    (pi0 == 8'h64) ? 8'h8C :
    (pi0 == 8'h65) ? 8'hBC :
    (pi0 == 8'h66) ? 8'hD3 :
    (pi0 == 8'h67) ? 8'h0A :
    (pi0 == 8'h68) ? 8'hF7 :
    (pi0 == 8'h69) ? 8'hE4 :
    (pi0 == 8'h6A) ? 8'h58 :
    (pi0 == 8'h6B) ? 8'h05 :
    (pi0 == 8'h6C) ? 8'hB8 :
    (pi0 == 8'h6D) ? 8'hB3 :
    (pi0 == 8'h6E) ? 8'h45 :
    (pi0 == 8'h6F) ? 8'h06 :
    (pi0 == 8'h70) ? 8'hD0 :
    (pi0 == 8'h71) ? 8'h2C :
    (pi0 == 8'h72) ? 8'h1E :
    (pi0 == 8'h73) ? 8'h8F :
    (pi0 == 8'h74) ? 8'hCA :
    (pi0 == 8'h75) ? 8'h3F :
    (pi0 == 8'h76) ? 8'h0F :
    (pi0 == 8'h77) ? 8'h02 :
    (pi0 == 8'h78) ? 8'hC1 :
    (pi0 == 8'h79) ? 8'hAF :
    (pi0 == 8'h7A) ? 8'hBD :
    (pi0 == 8'h7B) ? 8'h03 :
    (pi0 == 8'h7C) ? 8'h01 :
    (pi0 == 8'h7D) ? 8'h13 :
    (pi0 == 8'h7E) ? 8'h8A :
    (pi0 == 8'h7F) ? 8'h6B :
    (pi0 == 8'h80) ? 8'h3A :
    (pi0 == 8'h81) ? 8'h91 :
    (pi0 == 8'h82) ? 8'h11 :
    (pi0 == 8'h83) ? 8'h41 :
    (pi0 == 8'h84) ? 8'h4F :
    (pi0 == 8'h85) ? 8'h67 :
    (pi0 == 8'h86) ? 8'hDC :
    (pi0 == 8'h87) ? 8'hEA :
    (pi0 == 8'h88) ? 8'h97 :
    (pi0 == 8'h89) ? 8'hF2 :
    (pi0 == 8'h8A) ? 8'hCF :
    (pi0 == 8'h8B) ? 8'hCE :
    (pi0 == 8'h8C) ? 8'hF0 :
    (pi0 == 8'h8D) ? 8'hB4 :
    (pi0 == 8'h8E) ? 8'hE6 :
    (pi0 == 8'h8F) ? 8'h73 :
    (pi0 == 8'h90) ? 8'h96 :
    (pi0 == 8'h91) ? 8'hAC :
    (pi0 == 8'h92) ? 8'h74 :
    (pi0 == 8'h93) ? 8'h22 :
    (pi0 == 8'h94) ? 8'hE7 :
    (pi0 == 8'h95) ? 8'hAD :
    (pi0 == 8'h96) ? 8'h35 :
    (pi0 == 8'h97) ? 8'h85 :
    (pi0 == 8'h98) ? 8'hE2 :
    (pi0 == 8'h99) ? 8'hF9 :
    (pi0 == 8'h9A) ? 8'h37 :
    (pi0 == 8'h9B) ? 8'hE8 :
    (pi0 == 8'h9C) ? 8'h1C :
    (pi0 == 8'h9D) ? 8'h75 :
    (pi0 == 8'h9E) ? 8'hDF :
    (pi0 == 8'h9F) ? 8'h6E :
    (pi0 == 8'hA0) ? 8'h47 :
    (pi0 == 8'hA1) ? 8'hF1 :
    (pi0 == 8'hA2) ? 8'h1A :
    (pi0 == 8'hA3) ? 8'h71 :
    (pi0 == 8'hA4) ? 8'h1D :
    (pi0 == 8'hA5) ? 8'h29 :
    (pi0 == 8'hA6) ? 8'hC5 :
    (pi0 == 8'hA7) ? 8'h89 :
    (pi0 == 8'hA8) ? 8'h6F :
    (pi0 == 8'hA9) ? 8'hB7 :
    (pi0 == 8'hAA) ? 8'h62 :
    (pi0 == 8'hAB) ? 8'h0E :
    (pi0 == 8'hAC) ? 8'hAA :
    (pi0 == 8'hAD) ? 8'h18 :
    (pi0 == 8'hAE) ? 8'hBE :
    (pi0 == 8'hAF) ? 8'h1B :
    (pi0 == 8'hB0) ? 8'hFC :
    (pi0 == 8'hB1) ? 8'h56 :
    (pi0 == 8'hB2) ? 8'h3E :
    (pi0 == 8'hB3) ? 8'h4B :
    (pi0 == 8'hB4) ? 8'hC6 :
    (pi0 == 8'hB5) ? 8'hD2 :
    (pi0 == 8'hB6) ? 8'h79 :
    (pi0 == 8'hB7) ? 8'h20 :
    (pi0 == 8'hB8) ? 8'h9A :
    (pi0 == 8'hB9) ? 8'hDB :
    (pi0 == 8'hBA) ? 8'hC0 :
    (pi0 == 8'hBB) ? 8'hFE :
    (pi0 == 8'hBC) ? 8'h78 :
    (pi0 == 8'hBD) ? 8'hCD :
    (pi0 == 8'hBE) ? 8'h5A :
    (pi0 == 8'hBF) ? 8'hF4 :
    (pi0 == 8'hC0) ? 8'h1F :
    (pi0 == 8'hC1) ? 8'hDD :
    (pi0 == 8'hC2) ? 8'hA8 :
    (pi0 == 8'hC3) ? 8'h33 :
    (pi0 == 8'hC4) ? 8'h88 :
    (pi0 == 8'hC5) ? 8'h07 :
    (pi0 == 8'hC6) ? 8'hC7 :
    (pi0 == 8'hC7) ? 8'h31 :
    (pi0 == 8'hC8) ? 8'hB1 :
    (pi0 == 8'hC9) ? 8'h12 :
    (pi0 == 8'hCA) ? 8'h10 :
    (pi0 == 8'hCB) ? 8'h59 :
    (pi0 == 8'hCC) ? 8'h27 :
    (pi0 == 8'hCD) ? 8'h80 :
    (pi0 == 8'hCE) ? 8'hEC :
    (pi0 == 8'hCF) ? 8'h5F :
    (pi0 == 8'hD0) ? 8'h60 :
    (pi0 == 8'hD1) ? 8'h51 :
    (pi0 == 8'hD2) ? 8'h7F :
    (pi0 == 8'hD3) ? 8'hA9 :
    (pi0 == 8'hD4) ? 8'h19 :
    (pi0 == 8'hD5) ? 8'hB5 :
    (pi0 == 8'hD6) ? 8'h4A :
    (pi0 == 8'hD7) ? 8'h0D :
    (pi0 == 8'hD8) ? 8'h2D :
    (pi0 == 8'hD9) ? 8'hE5 :
    (pi0 == 8'hDA) ? 8'h7A :
    (pi0 == 8'hDB) ? 8'h9F :
    (pi0 == 8'hDC) ? 8'h93 :
    (pi0 == 8'hDD) ? 8'hC9 :
    (pi0 == 8'hDE) ? 8'h9C :
    (pi0 == 8'hDF) ? 8'hEF :
    (pi0 == 8'hE0) ? 8'hA0 :
    (pi0 == 8'hE1) ? 8'hE0 :
    (pi0 == 8'hE2) ? 8'h3B :
    (pi0 == 8'hE3) ? 8'h4D :
    (pi0 == 8'hE4) ? 8'hAE :
    (pi0 == 8'hE5) ? 8'h2A :
    (pi0 == 8'hE6) ? 8'hF5 :
    (pi0 == 8'hE7) ? 8'hB0 :
    (pi0 == 8'hE8) ? 8'hC8 :
    (pi0 == 8'hE9) ? 8'hEB :
    (pi0 == 8'hEA) ? 8'hBB :
    (pi0 == 8'hEB) ? 8'h3C :
    (pi0 == 8'hEC) ? 8'h83 :
    (pi0 == 8'hED) ? 8'h53 :
    (pi0 == 8'hEE) ? 8'h99 :
    (pi0 == 8'hEF) ? 8'h61 :
    (pi0 == 8'hF0) ? 8'h17 :
    (pi0 == 8'hF1) ? 8'h2B :
    (pi0 == 8'hF2) ? 8'h04 :
    (pi0 == 8'hF3) ? 8'h7E :
    (pi0 == 8'hF4) ? 8'hBA :
    (pi0 == 8'hF5) ? 8'h77 :
    (pi0 == 8'hF6) ? 8'hD6 :
    (pi0 == 8'hF7) ? 8'h26 :
    (pi0 == 8'hF8) ? 8'hE1 :
    (pi0 == 8'hF9) ? 8'h69 :
    (pi0 == 8'hFA) ? 8'h14 :
    (pi0 == 8'hFB) ? 8'h63 :
    (pi0 == 8'hFC) ? 8'h55 :
    (pi0 == 8'hFD) ? 8'h21 :
    (pi0 == 8'hFE) ? 8'h0C :
    8'h00;

endmodule
